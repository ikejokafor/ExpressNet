`ifndef	__CNN_LAYER_ACCEL_INTF__
`define	__CNN_LAYER_ACCEL_INTF__


interface cnn_layer_accel_intf

endinterface: cnn_layer_accel_intf


`endif