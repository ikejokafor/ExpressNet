`ifndef __CNL_SC2_VERIF_DEFS__
`define __CNL_SC2_VERIF_DEFS__


`define cnl_scX_DUTOutput       cnl_sc2_DUTOutput
`define cnl_scX_generator       cnl_sc2_generator
`define cnl_scX_monitor         cnl_sc2_monitor
`define cnl_scX_scoreboard      cnl_sc2_scoreboard
`define cnl_scX_agent           cnl_sc2_agent
`define cnl_scX_assertion       cnl_sc2_assertion
`define cnl_scX_driver          cnl_sc2_driver
`define cnl_scX_environment     cnl_sc2_environment

`define scX_DUTOutParams_t      sc2_DUTOutParams_t
`define scX_datum_t             sc2_datum_t
`define scX_genParams_t         sc2_genParams_tarams_t
`define scX_testParams_t        sc2_testParams_t
`define scX_monParams_t         sc2_monParams_t
`define scX_scoreParams_t       sc2_scoreParams_t
`define scX_agentParams_t       sc2_agentParams_t
`define scX_asrtParams_t        sc2_asrtParams_t
`define scX_drvParams_t         sc2_drvParams_t


`define scX_DUTOutParams        sc2_DUTOutParams
`define scX_datum               sc2_datum
`define scX_genParams           sc2_genParams_tarams
`define scX_testParams          sc2_testParams
`define scX_monParams           sc2_monParams
`define scX_scoreParams         sc2_scoreParams
`define scX_agentParams         sc2_agentParams
`define scX_asrtParams          sc2_asrtParams
`define scX_drvParams           sc2_drvParams
`define scX_query               sc2_query
`define scX_test                sc2_test
`define scX_sol                 sc2_sol


`endif
