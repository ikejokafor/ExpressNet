module dummy #(
    parameter r,
    parameter c,
    parameter p,
    parameter name,
    parameter idx,
    parameter wr_idx = 0,
    parameter rd_idx = 0
) (

);

endmodule
