library verilog;
use verilog.vl_types.all;
entity cnl_sc1_environment_sv_unit is
end cnl_sc1_environment_sv_unit;
