library verilog;
use verilog.vl_types.all;
entity blk_mem_gen_v8_3_5 is
    generic(
        C_CORENAME      : string  := "blk_mem_gen_v8_3_5";
        C_FAMILY        : string  := "virtex7";
        C_XDEVICEFAMILY : string  := "virtex7";
        C_ELABORATION_DIR: string  := "";
        C_INTERFACE_TYPE: integer := 0;
        C_USE_BRAM_BLOCK: integer := 0;
        C_CTRL_ECC_ALGO : string  := "NONE";
        C_ENABLE_32BIT_ADDRESS: integer := 0;
        C_AXI_TYPE      : integer := 0;
        C_AXI_SLAVE_TYPE: integer := 0;
        C_HAS_AXI_ID    : integer := 0;
        C_AXI_ID_WIDTH  : integer := 4;
        C_MEM_TYPE      : integer := 2;
        C_BYTE_SIZE     : integer := 9;
        C_ALGORITHM     : integer := 1;
        C_PRIM_TYPE     : integer := 3;
        C_LOAD_INIT_FILE: integer := 0;
        C_INIT_FILE_NAME: string  := "";
        C_INIT_FILE     : string  := "";
        C_USE_DEFAULT_DATA: integer := 0;
        C_DEFAULT_DATA  : string  := "0";
        C_HAS_RSTA      : integer := 0;
        C_RST_PRIORITY_A: string  := "CE";
        C_RSTRAM_A      : integer := 0;
        C_INITA_VAL     : string  := "0";
        C_HAS_ENA       : integer := 1;
        C_HAS_REGCEA    : integer := 0;
        C_USE_BYTE_WEA  : integer := 0;
        C_WEA_WIDTH     : integer := 1;
        C_WRITE_MODE_A  : string  := "WRITE_FIRST";
        C_WRITE_WIDTH_A : integer := 32;
        C_READ_WIDTH_A  : integer := 32;
        C_WRITE_DEPTH_A : integer := 64;
        C_READ_DEPTH_A  : integer := 64;
        C_ADDRA_WIDTH   : integer := 5;
        C_HAS_RSTB      : integer := 0;
        C_RST_PRIORITY_B: string  := "CE";
        C_RSTRAM_B      : integer := 0;
        C_INITB_VAL     : string  := "";
        C_HAS_ENB       : integer := 1;
        C_HAS_REGCEB    : integer := 0;
        C_USE_BYTE_WEB  : integer := 0;
        C_WEB_WIDTH     : integer := 1;
        C_WRITE_MODE_B  : string  := "WRITE_FIRST";
        C_WRITE_WIDTH_B : integer := 32;
        C_READ_WIDTH_B  : integer := 32;
        C_WRITE_DEPTH_B : integer := 64;
        C_READ_DEPTH_B  : integer := 64;
        C_ADDRB_WIDTH   : integer := 5;
        C_HAS_MEM_OUTPUT_REGS_A: integer := 0;
        C_HAS_MEM_OUTPUT_REGS_B: integer := 0;
        C_HAS_MUX_OUTPUT_REGS_A: integer := 0;
        C_HAS_MUX_OUTPUT_REGS_B: integer := 0;
        C_HAS_SOFTECC_INPUT_REGS_A: integer := 0;
        C_HAS_SOFTECC_OUTPUT_REGS_B: integer := 0;
        C_MUX_PIPELINE_STAGES: integer := 0;
        C_USE_SOFTECC   : integer := 0;
        C_USE_ECC       : integer := 0;
        C_EN_ECC_PIPE   : integer := 0;
        C_HAS_INJECTERR : integer := 0;
        C_SIM_COLLISION_CHECK: string  := "NONE";
        C_COMMON_CLK    : integer := 1;
        C_DISABLE_WARN_BHV_COLL: integer := 0;
        C_EN_SLEEP_PIN  : integer := 0;
        C_USE_URAM      : integer := 0;
        C_EN_RDADDRA_CHG: integer := 0;
        C_EN_RDADDRB_CHG: integer := 0;
        C_EN_DEEPSLEEP_PIN: integer := 0;
        C_EN_SHUTDOWN_PIN: integer := 0;
        C_EN_SAFETY_CKT : integer := 0;
        C_COUNT_36K_BRAM: string  := "";
        C_COUNT_18K_BRAM: string  := "";
        C_EST_POWER_SUMMARY: string  := "";
        C_DISABLE_WARN_BHV_RANGE: integer := 0
    );
    port(
        clka            : in     vl_logic;
        rsta            : in     vl_logic;
        ena             : in     vl_logic;
        regcea          : in     vl_logic;
        wea             : in     vl_logic_vector;
        addra           : in     vl_logic_vector;
        dina            : in     vl_logic_vector;
        douta           : out    vl_logic_vector;
        clkb            : in     vl_logic;
        rstb            : in     vl_logic;
        enb             : in     vl_logic;
        regceb          : in     vl_logic;
        web             : in     vl_logic_vector;
        addrb           : in     vl_logic_vector;
        dinb            : in     vl_logic_vector;
        doutb           : out    vl_logic_vector;
        injectsbiterr   : in     vl_logic;
        injectdbiterr   : in     vl_logic;
        sbiterr         : out    vl_logic;
        dbiterr         : out    vl_logic;
        rdaddrecc       : out    vl_logic_vector;
        eccpipece       : in     vl_logic;
        sleep           : in     vl_logic;
        deepsleep       : in     vl_logic;
        shutdown        : in     vl_logic;
        rsta_busy       : out    vl_logic;
        rstb_busy       : out    vl_logic;
        s_aclk          : in     vl_logic;
        s_aresetn       : in     vl_logic;
        s_axi_awid      : in     vl_logic_vector;
        s_axi_awaddr    : in     vl_logic_vector(31 downto 0);
        s_axi_awlen     : in     vl_logic_vector(7 downto 0);
        s_axi_awsize    : in     vl_logic_vector(2 downto 0);
        s_axi_awburst   : in     vl_logic_vector(1 downto 0);
        s_axi_awvalid   : in     vl_logic;
        s_axi_awready   : out    vl_logic;
        s_axi_wdata     : in     vl_logic_vector;
        s_axi_wstrb     : in     vl_logic_vector;
        s_axi_wlast     : in     vl_logic;
        s_axi_wvalid    : in     vl_logic;
        s_axi_wready    : out    vl_logic;
        s_axi_bid       : out    vl_logic_vector;
        s_axi_bresp     : out    vl_logic_vector(1 downto 0);
        s_axi_bvalid    : out    vl_logic;
        s_axi_bready    : in     vl_logic;
        s_axi_arid      : in     vl_logic_vector;
        s_axi_araddr    : in     vl_logic_vector(31 downto 0);
        s_axi_arlen     : in     vl_logic_vector(7 downto 0);
        s_axi_arsize    : in     vl_logic_vector(2 downto 0);
        s_axi_arburst   : in     vl_logic_vector(1 downto 0);
        s_axi_arvalid   : in     vl_logic;
        s_axi_arready   : out    vl_logic;
        s_axi_rid       : out    vl_logic_vector;
        s_axi_rdata     : out    vl_logic_vector;
        s_axi_rresp     : out    vl_logic_vector(1 downto 0);
        s_axi_rlast     : out    vl_logic;
        s_axi_rvalid    : out    vl_logic;
        s_axi_rready    : in     vl_logic;
        s_axi_injectsbiterr: in     vl_logic;
        s_axi_injectdbiterr: in     vl_logic;
        s_axi_sbiterr   : out    vl_logic;
        s_axi_dbiterr   : out    vl_logic;
        s_axi_rdaddrecc : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_CORENAME : constant is 1;
    attribute mti_svvh_generic_type of C_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of C_XDEVICEFAMILY : constant is 1;
    attribute mti_svvh_generic_type of C_ELABORATION_DIR : constant is 1;
    attribute mti_svvh_generic_type of C_INTERFACE_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_USE_BRAM_BLOCK : constant is 1;
    attribute mti_svvh_generic_type of C_CTRL_ECC_ALGO : constant is 1;
    attribute mti_svvh_generic_type of C_ENABLE_32BIT_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_AXI_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_AXI_SLAVE_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_AXI_ID : constant is 1;
    attribute mti_svvh_generic_type of C_AXI_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_MEM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_BYTE_SIZE : constant is 1;
    attribute mti_svvh_generic_type of C_ALGORITHM : constant is 1;
    attribute mti_svvh_generic_type of C_PRIM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_LOAD_INIT_FILE : constant is 1;
    attribute mti_svvh_generic_type of C_INIT_FILE_NAME : constant is 1;
    attribute mti_svvh_generic_type of C_INIT_FILE : constant is 1;
    attribute mti_svvh_generic_type of C_USE_DEFAULT_DATA : constant is 1;
    attribute mti_svvh_generic_type of C_DEFAULT_DATA : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RSTA : constant is 1;
    attribute mti_svvh_generic_type of C_RST_PRIORITY_A : constant is 1;
    attribute mti_svvh_generic_type of C_RSTRAM_A : constant is 1;
    attribute mti_svvh_generic_type of C_INITA_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ENA : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_REGCEA : constant is 1;
    attribute mti_svvh_generic_type of C_USE_BYTE_WEA : constant is 1;
    attribute mti_svvh_generic_type of C_WEA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_MODE_A : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_WIDTH_A : constant is 1;
    attribute mti_svvh_generic_type of C_READ_WIDTH_A : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_DEPTH_A : constant is 1;
    attribute mti_svvh_generic_type of C_READ_DEPTH_A : constant is 1;
    attribute mti_svvh_generic_type of C_ADDRA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RSTB : constant is 1;
    attribute mti_svvh_generic_type of C_RST_PRIORITY_B : constant is 1;
    attribute mti_svvh_generic_type of C_RSTRAM_B : constant is 1;
    attribute mti_svvh_generic_type of C_INITB_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ENB : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_REGCEB : constant is 1;
    attribute mti_svvh_generic_type of C_USE_BYTE_WEB : constant is 1;
    attribute mti_svvh_generic_type of C_WEB_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_MODE_B : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_WIDTH_B : constant is 1;
    attribute mti_svvh_generic_type of C_READ_WIDTH_B : constant is 1;
    attribute mti_svvh_generic_type of C_WRITE_DEPTH_B : constant is 1;
    attribute mti_svvh_generic_type of C_READ_DEPTH_B : constant is 1;
    attribute mti_svvh_generic_type of C_ADDRB_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_MEM_OUTPUT_REGS_A : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_MEM_OUTPUT_REGS_B : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_MUX_OUTPUT_REGS_A : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_MUX_OUTPUT_REGS_B : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SOFTECC_INPUT_REGS_A : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SOFTECC_OUTPUT_REGS_B : constant is 1;
    attribute mti_svvh_generic_type of C_MUX_PIPELINE_STAGES : constant is 1;
    attribute mti_svvh_generic_type of C_USE_SOFTECC : constant is 1;
    attribute mti_svvh_generic_type of C_USE_ECC : constant is 1;
    attribute mti_svvh_generic_type of C_EN_ECC_PIPE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_INJECTERR : constant is 1;
    attribute mti_svvh_generic_type of C_SIM_COLLISION_CHECK : constant is 1;
    attribute mti_svvh_generic_type of C_COMMON_CLK : constant is 1;
    attribute mti_svvh_generic_type of C_DISABLE_WARN_BHV_COLL : constant is 1;
    attribute mti_svvh_generic_type of C_EN_SLEEP_PIN : constant is 1;
    attribute mti_svvh_generic_type of C_USE_URAM : constant is 1;
    attribute mti_svvh_generic_type of C_EN_RDADDRA_CHG : constant is 1;
    attribute mti_svvh_generic_type of C_EN_RDADDRB_CHG : constant is 1;
    attribute mti_svvh_generic_type of C_EN_DEEPSLEEP_PIN : constant is 1;
    attribute mti_svvh_generic_type of C_EN_SHUTDOWN_PIN : constant is 1;
    attribute mti_svvh_generic_type of C_EN_SAFETY_CKT : constant is 1;
    attribute mti_svvh_generic_type of C_COUNT_36K_BRAM : constant is 1;
    attribute mti_svvh_generic_type of C_COUNT_18K_BRAM : constant is 1;
    attribute mti_svvh_generic_type of C_EST_POWER_SUMMARY : constant is 1;
    attribute mti_svvh_generic_type of C_DISABLE_WARN_BHV_RANGE : constant is 1;
end blk_mem_gen_v8_3_5;
