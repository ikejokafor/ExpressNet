`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2BUHvOFc2vGpCxhr2whtCiKPaW8g+8+86qUuUvEkmbF7gu+Y/R2kGukxTchD16S9
2laKr7HC1ygyziKpqHWMuDw6lx/XiuKkV5Fzz2MuUVyGSq8jI/wqguaEux5C3HM5
U58K8F0NNOjR8wDdnD6RivuEpjS3VDwWYRCyamk2hu9WrlCxuOMR5t+aJ7Ilwq3q
kRwtbGvfuHlwrE2M+qYh94ArbXa8Xk5C1izsDwTcXwoKqbpIfGHr3tf+CU/oblQh
b/zUCwLffZkqzzmwBEjRQMPS0LgerbsC3r3RKcr4Md35gTHBA6V3qOKBtapw/JyO
ibAcQxIDBeL0XqMR4ezZKxI+V12qq59QFrTtRXLkNouC3rN6xmd4jaUwAq6zn9q2
8cXIZdZHrCQc+nfrbH6Za6jF48W2FkN44mY1IXTD27DiMCUCUe3S1BEBukefkJ4f
a637ref+BEzD1C+rQyfWFTBmSqXOgmTiCUfbhVr6xtUy8KCAL1zu+3/3S0rkp7Zd
zXYlgQsuI7DpXJzwBpZeHgMOOHgJCtCkFFk9X7j+03Mtinjezx7z0h7nmEVqe3Uk
m0xyDqrE+ExQKgiDJVDBdctWbLPLKRGBqtRPC/Jk21lk29jC5GvJyXgafVKJMttN
orRGgSfkC5roS2uYKT2FEQrDWCNDnEfRFKrFYLehGqYvEhujbMfx+8I5sn1qWRc5
+3qdCQA7nPDWCSOo5xMoNZCAdCvpYqKs2k2Hbr4z+AFuABeZDANbjES6QTtrRmDy
VY1/5j9J1iCjG7FB4xr040PQu4pz6IP1vJkNLk6AYv1khKQzhNi4TQIz2HYFrzx/
J1lqujUGY1ylxBCr5yc6p4AZxMVXTlevVK8YdVcZz96chu+biAwnWYdRZ1bSE3IL
ooyJwXhaUDZr3Flpy1DxEd92UITJp6+dPFA4W29MyvKmymQbaqhdQ3wF8yz+Dr61
U5gg20/TGh3PyOuMlYlw7CEEGemPQuaFNMyxQ+iB7gOwQ5zHhAQlhI1BAjV9IKpf
5bh5clc0anMUTmJGsRM9IwFN5qed7/NHK82gZX52p3/CmMunW/FnhrSon/Fnzn5N
mqNeVDqAQHQSFdmHCLA0QMA/43Y+azlTUhF+ERME4pcrUsJcajfv+TdVdOWF8aKW
pikqWRzDFqJAREEgGWMdJ0RnUGBtTrSUBLaVzUCrjWuHJlKESaMANETmWqgIo40U
huxmW3IjvG/7W9NnO9C05qmLAST50TKiarjEfXT2Nh4OjjveXvafZ4vAPYJSlssk
j7i4jeJkTNTBn9pvATvLcbCS9R2sPH9UcrxcIZWDzKzOh6HR7q+4DOdvBFfAHHRJ
Y+Mx3SJwRyvkJ7JInTxQsvCQ0Bv1b/Ms/NvI0OFT3Yt46Ful1K7ZCQYZ/Sa5y9rQ
9k+jW3sr5/+xUmTspuuqiHAzfzNmZH+NAHEc9ZZ/h/44ILxZ1/qnPeU0yXgmRvhL
ECiOERUHShJNx/N/pXi87hew4LfFOpC1wwV1bDLMSv8fyNscXCgglqu9VYGZGKmK
4VlKLGJ6OVn+y3sGOEaKtSA2rnzk1RYSl57EaOa4RvE18BA9nS9MJOTHtlGvp9iF
bv3BMIL3GScSSe/+cxipluh0cC86B+7aS+xGqP113sS8kXg+KpYyV5UBb/uXkjEn
4hF++P8+8j3HMIMA38sCyMcs7cXeffsrz8eDODjFXVj4YqotKXGUKwXhMgaN0+e1
HUn/iDigPik3a9m1C4ABeFoi1QPwMA6n95iCK5nfrOeJPSMaSxRlJZHht5bSmny+
SJaJ652CV9yXHxu9h+UdzBVa/zlhcwlLK6LpavaTMBhtlbdxYoKzEMSZR47pgi4i
/mObnbZDqvrP0ac5tRdZleobV68PnDMHD0iLPyd60dxaY/WRdjJHeCGsStAQ1N/Q
jK2aJXT6Gu3AW1SKX2VeRdYdK+GM6srOO86S6Wtiyr18klp+sUfyz55mnokZauaV
1bY8z3aIoHz5Xi1PH9lO2B9pgIx1nUhrhRzXD8S12CGQeftFm29KQ5fdmSdn2zDa
lcRctVQau+n8yyMja5Q1jLuyY4kwdlMrwmnNrAFoNMGN3tPRXWbSqu3ZM8yaCYgn
tE+AZUPEh0+H627cL5oPlqtYS6FQfuj6tkdVExg6aZCWSAlwbGpnfsDosKBDQZNz
UYQrgNftx/s33JTWZYz7y+md4/CUCMjpIDyiVZ5hbjGh0h8D4/ANTguABCk7SOrc
ahMIDfPgDPpF42Ax7UUGmMzCqLl11tjZZAO2e2LQkgoxA0C8tixxs4lG6oxlXY2t
RYQKAxyrwmKLVB2sAE20X17zZ3ikYcrDNNJCVGUCXKe0FvX8Qk9DYcjN4/qWguUG
oU83BuRzT82czTJBTWwfOsXrL9EAWLkVLKxz6C0XcKRs2ZVmx78xHsAY+caRhO2U
vy9eAM8BWsZMalzsad78hd5kQOOWlPRS8dKGZAecr4KqRnbwGXeEu1D9gQ0qLLB1
dTsl4fITYAUJDp6Qa2/tvMcN5OLpDgugAhQnlifyczVE9l6Vgt780Ap1QTGCV9fA
WdWAbusd0G2ovwQNFyLvdih82Du0+XFDj25vz5c0GuriXfxB3htn0JeAUW0uqFLQ
QYqdrrh+ru6jNGF76AnxuIh0wjMLlAIO4L77yIrrAoa/P+cer2Mt7XDuJb6G0bqK
TQaUSwMAYIcyASJtcu67ETNWzPw8On/Ak1TttHU+VJzxrq1cfqgaVsgx5QqY0zk3
+9iTYIxB3eralq2OTyBb0+AYM7NMtZxwSCI1jZkpu3vz3KFE7YAlczxrx8xKabGX
8/oFYZxQU5xQF+ho4fOAE4+6TiiLtSjDSL7BbqwLOiuSrEjo1qivb/WVzjKvUF5/
NxBvATpZGNTdm1mnwL8xoHYS9QRmMBvacABwrtkIUE539M5UdzWbYHgM59RMcF33
2nkMU3TGFZAYBCtPi5dmwh3y5j1zzbQa0ZQRHMUkkpsb9LcPxldGk2M4GVn88Aw9
lhAYh4NYr1VLGgCong/vny7v2usOUfrWu96v+ZkH+X3d3S5NBqxI63iJyI3v5gYH
OrRH0WI4iMM43en0NO5ad0hgXsllu7S+NnDV6qPt5c2wTndl8xWGTl30zSzh8Xup
cQ9mfTb9b79ohC0q8Qc0iU0uVjyDiO9CGxOV0FhVjKLj1rS/BSNe5JH0YF1CKvN3
OcyViCjtf8KijEJVRdgDe51NUzt8sj6+Irxgvfa3vaUkQ3+HsLaa6rAplUzXxE1E
iDyh9ziEJpUfJxkKnGpq5QQVioZxQbwIExp1hxAIjVOviK52/XCLRqStTck3AvFF
m9Unfs/ad4F5fGcdM4FEHtVO0St8Nk1U0qSJ3dgJpvTUVVM811rNI1629qtVB/6g
mS/8qLQ0YlC2CWkSHVVTSFWKSTW1eUz3YcYyn3UwQBW+oRVwOK+zIXF6w9lgTc0F
gNrzq7872Ig8BnWCyJjYkJi6+C0v8Rep/AcdRCVijdirCS4kOIh/Bmp1a6r46Qj+
OEriGEC/zoksxorGRpLeB+NO39oiqFOy4aN1slMRYfcxVYuvpTsJMKyeuOW0KgLc
DX/oKh5pZURTbJWO/7u7xwXMYCyXjVeh3MQpTEN2oM8PSGnQtl0UwFbeU87ZyheH
sLDzr88Dc4lkMzo7eUlq9Dg2rZcErHiZDdSPYC+TSF641/V2LqF+xPnMl2XmY7bm
CHuRTMtEUJYHR72c7CC8KhD2jgo2J7XmaPgCKvfTzGLmcMhCuM6SBLY95UkxTNT+
ldFggo5fIZYzHb+B7n+yvO4HIcWwhUGXs+VDxCwHY26aw61nUAgtkxgAOoBCm3t2
O3A61fX1FbsMPH9TCiaSS2+fE9RPBhJp+08vqC+q1/b5TSOclmtzbZsR7ahwBq/j
2mTsTaDX02WYSBlwygwgTVQIRkavepuUtXSSNDbUnxPkJwHgfaBJtZgk7yiTMiw4
04i3uylrfKoE8HQU/71bCafWlUe5f4cHod871Ke5vCZ0uTwtAQdoIwRzUVkuj5tL
mJgHaZq4Snr1RdF3D7t1AwF4dIxbm7xIfKA70xvQ/cNb9HlxQt2WNBe8dfUZ1CCL
sUiV047o1hDtxyJyM87/VcwB+AnguSXtaFg2Lq+ZC9u85D+G3axY1WMYK4WT7V0s
mKaBoEWxeCAoilROdwTI6fKYjGnktBOqLxBuBAR1nlPETX00TswOKluw9b9lu/7h
DGA4wdBZN0Pa3YV6vJyf+yyeiD7e3QCG/NC0o0FuhmyCrbfd3NlbgQc98pOCI+rF
/jull5Da/+qmE7e7+Bwk8fRjkh2Pzcf5pMnbA7rYQ2doeM9A8gn03xFbrOPdlLJA
5dJodncSQASMLsvgcv7+8xmHiDOIpN5gkfJg2hSxea8CoIPMt+wugROX7bNb04KW
QJOT/U2VnYaOhvQMNzBn/FVRaeMdjzI/QFbzpSHh92e9q9W0ArZs7JjVZ19mUsL4
BnHS96I+EQfGvt30K5T2xmzn4q7NDL2Dz4ssvd7Aqz0JInmsMtDrj3Y8HqJpf8Y8
sl9hDR+kAqo91BgDAKdQjZn8GVyvxRB4RYAI10I8whre9adolQyat0pz6F3vIh5L
ZgxlbuqEXvJ6/tN4QNbaUMq0XMQHQVOm5U7Ti9lLYmNYkF4x/EBasPqHW0DWKxQS
wjZ+XLv1FYpFD1PlodFceRXaH7HGQMZm9+l5oeqLq85xGhSVrEZKC5wxAIDTwrbY
4X0FiUv7nN0KuB4IVZfXFy3WwKikS4WVjKBMMu8IF7PzBTF3rWF034m0mBR83ZTR
IuNwK0JRxjxVJEsCLrBsP40E6rX4SVWGSW4xpKIkTr5UGq6N1LbOCeMiD0867ucE
D8l2tKrDn0U4dWSt2ZkPydXJHD2Nd6XmaSKpBM2oFT70Fk2dS6tCHDEZ1wzQNLUU
M1wtUs3yzvvxjNtSolzRHoHnVJVSxr05VbelEuNVQOzoMaqKcUxykBYTNYNB3nUJ
7bv+UmLviUZEC4yHCEqQqz4kPhbY7lnVDNZjHYl+obK4iRc4lLQ+BotnUoo3zRpF
2PkG/AWY8hTcAg2uRXhxfDoi2umFAbA3YkZp7+4kbmadoQ0HrWkwu1NZGGE7RMkk
mJ0B6wHb2BfCagHBp04exsy8ChooKke3qEx7xHjBu4v6hMM4fust5CIS9jipYhS0
yWXLJepXykLcK119j9iqnkEMPX2DaIXqQbphl7s+6nDlGpShMPxxzz3TmQjHte5J
L9C8LXaGuN03J2EAvRj9WXdGGxkQMTGmAIRHQiOmuPSFsF4P6r0xlgvrtndKbnmn
1tMHw7oB7iOflLL2pJjtJJGOq8zQFAGRFDRhUjGw1blnEVxlsxYsuwl3V67dM/+q
m76ijLvICgVgqxmNEP+F/K1airOqFz02BuVNLpUgAmNp3noF5G6NoEPvPXY9lj37
zBKYeLAMbLbr8JF7AiRmMRoGARiwwSfKbBh4IFUcSNcE/euSSyanVPOtHPAdi+M9
MYu85vMCyW+O0SDXoD7PBrfDIu/OCXVYjlF7xVc7obBrZxaPqE7BF7Y5htmDs9K/
xI6jH8IdsJXdSPmNMwI63flB0ypvYoV008sO25BAVmx6D6FnvivyjI3C01Lkkt/I
QoTkmAMS/4Tk5fwetCi4r1hfn7VCahK5465280cxBZhO2atI9LirKeq635gmEVCg
brOVpavwLwpgkO/pw9eAj1tukGTLBqlQI2C03Wg4Aq5q1B/hn3jU9BmfyXE0qZmu
cOdARWB5nVVvPGX3+q/lkyWt+UWFXE7lB71YwiO2q6Sx7ulW2a3AWuAj+2smYWW5
SjwJ0UvkWUeMAQlv7SMypKhnpjs/3MHTy7SejbcEdOfTzEAoz3H4SUJdmf0dN3Kc
VRc8XQ5gUMrZXvvCNdjk2JEwhCIe1cbgFgGUFR3FcsoWc5tEujnuuZN6rMTsw70H
sMLzJKAmzaqSPhuXp+Grg+M37nCUb8ShhWrOBVa+waR89Uq5jINEtlUx0lCngxpa
ngtGi5uA42BHm/KsknlsqM+GGBIRwP5mNGSjcGVQI0ubi0C/7fHZJDiJM7xVd2qK
TjS7xin35t8IihTuf6q17p56i8kih2KEq3Fe98mL7CqJ9ovfytuB7xr//esdegKf
eWg3Ug1cAD2C5u/RevSB6CkjRyjyQt9ktOb5kArCg0KoFyS4y9b7QShze0rwzT8J
rsm6uHN0G0pjwSHYG+CcNDh/nSO73mOmSW84nma6pUhRlav+hq8eEM6n0pIPo2oT
cl9MNWx+XEwMJIciHyhj+Uu2mRwn8DdJ1Q63pfBoWGO6S7ojVoZFGgBV8ko0dUhJ
RIoHdeIzH+Z5GukAnm9yfLJ2/x4lLNuV77LC8xtsLIE3xRAQIg1qY1Iw8sHrztWd
RXrGD5hoq2qzA9iituHX3h6wjT7oyQvb4aE7za9lrrFGNW0FqpV/mRSdV033C/Ca
BFtC4uxcytoq+wCLt0qXcK1sXhHmJMV99LJxPYKAVl63hUo1cJg4LHJN0URzZyF4
tkUIGktCsHceTr9BkKh6LWxoAAa4Ou1iniJnznNERVbJcgjwt6YcyIdOxUDu6ELI
k/RViVNloNfmVPepF0/bFTpa4joeHJ90gUClxmGtj27z/MMTagli/y+kHolfTBSz
J/OPeQ/XSabF6pJPCmddM88a/bDzcyCmU6VWMMXE8F1fMKHjhz27b4UHBOai4/M0
63Rd4zxcABILb5yto9o762lFB6PcPTYmzmVqqpJORA6Pz584uZyn0D4O44I4+7V1
0p26ms8bBznWbhupNmQKrcxo+iiXAatKNcG2Ukq7ryVSoCT521VGYicgnQUU76d6
ykNH6sG4D/6rUz+KAGpNK5oiSYtBF9Sy7iGl+iY71xqJ3CZzMpFvkmwvXMtL6ddY
thtiAYwK6TCC9N6AUcWwtJh/4QxLj5wFuwPvK7ggXBBQRi/UVwcTWDGcrhB4EaBr
qKh1J5VM5RlQZx3VKzgPo1AXwPhMlnNYkWB/d2+oW9uaOBE/kb6uI33QJpQuQQ7p
wBvVjVC9tlzwg0IuBovQj9kUeTfqUFyukvOM8xa0H6pSZUzi/NhePov5jhjGkNzD
AiU7KD2PWBtMEM0sBZIaBDPSjAgM9EQwnbIkn4ai8oX9QAgV51+PKXdnmwfT2xvA
IZVIyruLrPXJ6zBtmfb2IeLZ0Q3B58WqBwmL3ahcNv6kuLFytwMt13LFfjYn5NHB
eNLo9UdkAJ7p1ePdnsSOilXgVP+PRhXCqWfnhRh19+t0KG6tpA6ckPWirhmUiBcs
dMswG/eQSYOQdGIDQcLdQmhcreXOAiuGCnSL1l+xN2zmFs6VL7Ty2QZHZ9Vs0dTt
rA7vAP/jy88gN9zU4yVUE8Qud7qaYk+op+jbT9Z56buvckEmtymM5F6dAvJ0pMD/
TrvRzBTE0XNuQp/QGFYY9Wlfwl3on5jnyXbgiPVTbBpq7jcwYm/U62ami9dC08oI
xJg6RUbp5tmrcG98DBnnX/WIKJzKHgm2F5TcjxDlPc4//hfbXNuE7H3kPGHlvePX
4XhcHaS+NFApBvCT8i9hAGhleDpHoOWxx3j85En5fiNmeWLKh8z+S/L+Sh74pXmf
nq3dzN4v7QkdnSO4vCS3JA3Vme/7DWgYAl+jWN4fYhuZguVoRjmYigN45L9mBfoQ
6axG3rzOr+yE3sOrVd1SliO7Qg5Ij7gg8ZEVtOmYvv/OZtbzWw1aOU9lg/y8tjKh
r8vEX7pLFre9OdNFPAo2QXmTUMZnt2O+5KmHey/4N+Ar8pVCPGtkMv1L5NWI8XIJ
OAUZkHVPtxNfjF55o+Gmp38+4luSqp9yWAxbGtHZCjzMnCXRJQ8Qs8pxtdzohJZz
aeH2xRA1A2tgtC7EpyZ/5GUsahnVCZP1Immt3Mbn2Uqlw7SvWQFRJA0PN5Zwn4vB
teDywcA7DYGzXHB1S6H0aSI/6nzZ5PRyHXduRO9/oX3sFqHt+eBY6+SDBq7uuDP6
KPE+THnWbdj3Rwt4pKHHDNg3MR5v3yEWFOi/+rrfrYV9/J/OhyasqZHLgwR0QUsm
rUsNdUo8dKvjEJxtZEOO1vB5UBUpSmr4U5iUXa412J6y0qOly85mdZhurk6iufrv
hgyhQd6IhGlkcfbu7H4tvAfgnPd/oNI8Z+UPv/I7XO1gRc502MNSkBIgXjNgma+P
wFur1vvawIB/NfBwoqEWJUYohPnhce6wjZ58kOLMQCa2ggGSSpK3oy6e9BD1i80/
wY58oHm8WGrUgk105P96UsKIYuCN70oHpFxD6AJdeOz/5cNv9vIy9LqHXdqJuKTc
bGRoA2JvJ7E8V8GAv9nOgR/ts2298S21As340cu5JmXMzvkL2x5XYhzQ5pm0eY1S
c2KhmDw7pXAEssH+E0hQGLukG5LN960nSTk/b7VQEYhty3bDyLOp0fpQp4y0+cPV
YBGIqyyAT+T14Kn7v8NE2IG4QjRDhxc94nJ9aG/Pe3jvtZwWYftyj2hGnmC+RolK
7oWPeF81CHulsJSIIZSPbtq8z4rEUuSXt35omjCqqgKgEQ7ngcZbxQLi3AXNUGx7
EJc5OvUqiKckewq55+XsOvVDshu1pDL7ph5DOJuofjGnSPcxXexFKASqMX3JdSuR
l/8b5tcxzeJPFzmO6/FT15acViRr8pE6pQS7TmvOuxVhK53W479q3KHfY3+RU1v5
2Ud9sAn1sw5oCXpZZQBilCh9s742v5byxOfV1/fHZ2ufTgR7e4mNwyOUG4ip6mZ8
fxl7Zji/nnOy/N/I8K3atxqMv3Sg7svQ7SYzRzZ5lIRGnx9GYwQiWFydvV+wNQqS
0cbcx6tE5Ha9thFGqwlvtaSMoNT6MfHnknGcDj8lXzFDrplorW97ogqRRH6fnnjH
CrjXKDFIowKOtObsHG+dMPbILfimEYrjmdZK6AxHAjGwAvyW394KC/BZXvtsPrD+
SBISKSn/11Pp8P1shWKu1uLYp4zN9Q07p1AMRb7nKEPxH5t/WN1SV35g9G44u7Kf
MLpA0qnKBzqpgZip6VPUFLa2nplS1g4x53vwScA9As6gw09q1vezbgCv4+ObgePs
O7OG/s3zAgQmtm8tUKif2JyYVChlbjbVM5F7p5usKfIbFuKRKKnNSDsO23KAVxn7
/lI0OPPFnjnEZRWudXZ3oGJ/84Ke5uQyGdb89OTFbF5qPueS1j2CL4Vf8+J0rh6D
eR4qps1YYJp6GhmbVQ5fcEYPY1jGWSluzjZ4LuxOHghTrFdrwzhZeEExfhLqzdBr
kEoL3qHnMs8uOxEtWBxU7c5NtPzeruT0A7TdXqLvy9JtcsxaZYeFQia8GOMzvDXJ
Oc+PLqOeBv6Hm2xmyHg4gP/n+F0i67Zvi1sTuq24LnwhRV78EdrYxhiYwcgm3OVK
+8p2ozqyRg2NAZYMv7QWSi21Z+GcbmhLc5oNKA49lHm1hkKaYpQFhFBmK+GkQAv3
WZinIZp6QoluIlJKcd1HDScplU3a1xn4oR5OuinPD5/omR5Nw0z1TX0NwMzLCZVD
cF03P5vwYRenlyq5y6S+6OI/i6KcAwhgyfee5DKCqR0MLv1nJYYRTdGJZntga/yU
v/7oApsUZR9pxvseceD7B5DgyzhzN3JDfz3sTfEnXZy5a97wu3mVEEW69G7BkyoA
pdQqweefZ+C/nxI7MCf8kq5LJOnRGtXLdFoCbr7f9mmzmhT6JatQ+wHGLEmjzAnr
ABXM5mqSm8Mf9y4xEwJeTFl7WOrQQSjAWOqcTL/LLjZ2F2xZQ9ZQ9b76ZqYi1ciY
TEq5nGgo+zr7vG0K3lhZkOgWXf8GL9x3mGgwjRRDf0r8+FYHYNVPZU9WtjwL/SwV
2+IeJs8dYUpSUskFTcFUDagsUaM7/cQ0u2j4Qqw3CE7kaWneduyAgG3xHgfo598M
6tZ1SRzdjoPALZfsHGk/hUBumLtAK48LqBOtCB+W8pPvffEF6CPE6O8vzhrbEAD6
HKbuxXxFiD8agX+1vlZDe0gYw3mASfdaxY0PXsG4x+N1vqQ8W8Hrj0N9C+pnCbZL
qMZHITgFZDpQbamfpOVCKekGTIxbfLUM0f543XPO8Db0JSGqyhSg47vDMI7nyniD
wXXS8iwyGDmhLspY5EGIU734+kfxx+PAcbgUl4VenbY5WsF5RJOXg6JJ50C4n5dX
TEEdOVIjJ8wQCkuQ01N97XMr2y95HIyZYblfhsOC+5Qe7oJ2EIxNeufhIgFFmQYd
mqD+OHpjAqguwYjdZhgRHBdPmcc+j71QcGWpSQuNVX/MB+cO93JnmKUhwZ33fFNt
DeMPkYkHYvtFdPDsmVScLK39J1ZsdCokrSDI/zRJFQVHlj7s7weSsQk2Nrp14+z3
5GUN0SFXqYmUvLpLjTo0mSMIbODusidB32Ai/fyrITjL/70SX0F5NzclzlvOZWpd
jqGb+tGgOxQMOFdK59CITg+C7A0tJkgvXatCQwKauQreVW3kTajSOp0NtEyTlZ6d
fjgPlCBcaKcTUuo1k2gpv8hSHuP4rivqKV1OxY+HorVibX9wQBr0thTKklk2bS7U
nrgysa3amc6nY6XLvS95SmF0WVoqZ0lx3bqt9GwvH/iZg95BPohgafV0gtI6ftnT
5HhYKgtUoa1cJ7PiqlyArrKdwvMKlAHdbCg0X8Ognt3Dgk40cNqNm0R4IB6bYuiv
kRZpiV9qImhXR06IyOnaie7liR1184fvBnFuW/isXGZPSmw7a006GBpo6bFstdsf
5jXmgeWfGM5d7H+uAyypgKxmwlE4NrZuCxD/f01BgKY4bHj+nkjY+NTZkG7OIjc9
0dk8V2d98hkGz/MAfYez8H1po1ME8J7glJ1T/2HxrUyBljN+P14qXzZ0+XCRi/yR
tTF0b6+SgUAiJhmtEQfthQqIrdZ6yoIhNwho86xfIzmSQxbB/ypBrjbObxpD8YHQ
5WzvExvZXEWTUPz5mVjLduMtKKDVSqO2O+Y5IHf0ov+S5zpXywphKly6thWEMhsC
NYs6PxQqUKZOuzJH1pyfOPbbQe7zHnC3SfFD6fHPBSChpc6WFTk0IbDJKS5wzlF7
ZWSGgwRBlb44IaFytVzYZj0y2QP4B0yQGVO17bAmt4iaHboEzG21DqRPR6p/3+gO
leqsG6KHbtgvsDj1g2OHM4W3bpBh8rWXcib9qFYgUTx8iaMuNfGP6MqHQlPqnKGL
kMEbQvfOY7MUju/W/q2OUJuMYn/xRZ1zz10dSfeK4f+mS0R5XlOgMQi7X+VvAbF3
wKoj3pHwlU0ceqKRJsCsTmRo/g3I6QZpyM4dyOGwx+Due8OcyTdjK/HqAvteEbVn
sPfIS8KlGCdPkH/yE+CgFqtPfuYp8edSb3FwU8Tdqu2HjeVSAp7GDwqucIgMo1r5
rJnPn7xpUDrAvF/LYQFzSU9z3SL+NejjXj+uXKZB8n7En6xKvqHs02mXgyz6RN1s
9z9LIeYD3VVeQ/nM+7CpjBosNDMXCOPU7Z8Hxke+NKs2BsbFsMfCogyqORAnf1Eh
jrvi7Xize/Phs+v+MYGVilfwvzzjIPwCCySRaj113EwKztg2I1ClxMw3UxjfPjGt
5f0pId8Dkx+sXe4LCTHOU3FfU0imUlDORrLf0+M9TpPCQ/NHDf33M2mv4gdvWiRW
abvZmHNE2YPNxs0z/P4XEOtG1LDvwxbfIaJz9tWkWdLtWBcAtDRQ7DbCqPeB62td
oTFYz7pmdUAOkJ7FSsuvtXUS6Bi7c+PwJTI9PsAF6eEf6ZZlWr4d1XSfbGYwChhS
97XlfAf0E+YZ9VYefHH18JvuHlNHkqWUUDAb/8NtbooIeVGuzMKeTU3Xeq3pJkNk
lcoemig8MkdYlpZ08vscF/AE3d7k+eA2uJ/o+4m7jwGIWBVlN2q0sqFtPwu2dePN
W+YNwknRLGN46i+Gn5oJQb18mZF5pUK2p00FzQ0fi7UenpvoyLOxG5nU8EY33/vk
rCkoJ+m6jPCHG1Dbo/Pyy3/Y1kca23WeTRglvtp+u9Kf5aUxa2W5a9tFNzXzFeNQ
61LU0jaApcNF/iKllD26/PvJo1zjtfomVy+Gm3ELOgszg8YZaYQUIAJG6lUOVg9m
dwB0kjK6M4GK/3R4zffDK4WVMVG+Pe5+G2BPnTxGa9jCvWzy4wIrbtgz7xfp+3wC
vn3WM94MdSGwveGQe8xmsRY6vGKjsxbUvl7QNxvnawniV/j2tGolvf0/AdSsDeqY
O9fWs+P2t2kyqN9njYIqQ/1mf1nIR2qO+0QOtheozfk/fkK8ENmwt89TbDw5wLQ5
yZsnsT53//pzA0UWIGWDunVWtdrBfYds5KJqWo/S7OpquZYEk36ShvC115t90kM9
+hDcj1pk0St/NkLv9+76HHeB/U9QRde3SELX/wTKqhd1rJ+Z2RIyGXSLev693kyA
Q98DUSJdYi/1nQGpwayAbDQOFa08IkKzLMyl24aJ0UE5D5eNwJR77vya4fS+dTzk
2mGjuN1VtM58E2kuN71ixDnpT9kUuvJLd7nzVDG5mGp83J4eH4dxw+9UdsBEc+gB
y2I1RkNz2fG50+702LwH6Oa7zAeQ4AiJ3uv1sPw/i7dMKkoLAbefRm1sETXEMPvH
T6JKbHL4RN5v+KAKdCG7ItOb58yo/Yqp/mPrgW4dKlVI8FlaTh4Tk+8nqy7r+wRy
QjDrYR/tKuRZkefXoN83gfJOUfXqqG780HUkFLivg+oRoML2lvIMsclDterg4M00
CeChXuh6p6NGfCIQpBbiVZ8GHIKUvyNhdtBtPEUpV1j0VTYS+BVbhUyaNIdRjfy5
lW46jroXEJVkC3LYLWbrnWFvekxtZlyLNn0qrTVUW0zraMVrPBa0xqoy6BKJie5t
jo5Ausyz2VSGME60Xd9sPo70apzLKCAhMmiJWOLPpGpiGQnGYK2V5V3usPab65+E
GxFVGBS3NcknC/sNwH6K6gQiiVjsiYE+nPTSMbGn2gLJGqd2K/C4nVd/cXg79h24
sEdVc8S+up5gSfcGHxMYuLbnJZ3BdAE49YYKZFja8pqQqHo/tpwQE5eXI7/2mFoX
8xvvrG/bVuslE3ZTSRQmlPKDBfJ0FWXS3Q9dVIPHn1w7GS0FEnfxZTknbIBkK0z0
oguagxNHzR/mTD1ZlZwHMkPyu0wsDGlBonQWYSyUecbINU6A3/ja548jmd6K5vfd
1HDlNKD4JdG76zbYiVDIaWNnvZmHhhYBMnW6/wms/BJoJ3Y2bq4mf3fXuZLnLxLg
vvNONLbcHYRTKV6oBNmTER3ZrKxYtjvsJi9bKBhO7ER0lTdUgrseqRFKgJcVnfnD
gb/ldN6i1JqEf+p6v1RRD23uUTahqp2OxI5dcJo7ISRHLQmDWepCz6u/3WX5zbyY
d/Yv7Ovr9mkJ5bdVCqfuaHqsues0n9Kcz1dX9zp8tUAM86hliLaD+oiKr7wKcZAG
KZDlP3BTapPFm/GUMsuTPNDvnb9fyADEBjR0mQf3r9n40WlOtpigp9LanuulTBu9
CfDg3j8xc033RqhT/YJaWsmJD2U9z9jJaFXb7qSeoLDo+/qSOx8CKo3TCtzEhASk
6uWtBnbETJjCYZ8P8pNsB+5m4UPApcJZ8LNqsAIiZx35bga3ZjViFjKZKGa9qEBQ
MmJl3IQJ7dl5VdNxBmOp3kYmIv5CXUBE0lakb9rVawrlo5vTA4j5mjC67IFLei1G
kobDTEEDKSwPEwLY+hxK3/6OFrx8mvoZH0jWoDR+WwEo/7ykyXJ+b+wMLxStcTml
9Y4My5DANgRo0ss8zFzJvg9n64xIx50irtg/32Ny/Zri9oOBSpp6Jx5FSwHax0w8
1OqWvHXaS2M82A65MUkwS+55jo4a271wyTJr9rv9iZFo3JGJ4Uv2AN/+KSLmrWNF
l9DTEtxRSqRddHmvBhqxpLdK3n/hU4l+bBD2VrANOrICoiZL6rVamBeV9k5q9pB5
/f5eM0kgPIytan1WLcDMhHwe0gx9u6V9pDEoL3kujCeK/xJeksgIJauA2fcwff4E
XUsjF3VCdd2yfpivINU/fkFX1o90K+lvb6IHBOtOIpfHpq4L1Kz9KcMQgJdt1ESi
z/MCG5PPRSdCJfpt15ri/k2cjVc3uiWs79hHwfcNYQ38XhhTdvBoELzQtj241qU9
Yyu3ny4G2Obbtd2eRmTfq4kvKrNcWrpIfGf8+tPez5ZuYtAYjOcFv5kDhdMCLWK0
Y2P4UN7j/GXq7tE4QOJJSLAsLJx1bEpCtgAMbE6urcIakPetBhuGUoImAkdaPyPZ
VXaLzBBDJ3RpiEFN9UKhtZUb20yQo27QqDJUcz3wZOJvlh9NTVvn5nEj5KDHWsbp
B5sMcAR5lmWIo5BogkqXZv/q0tJ25T1xcFHj9LMrI3rJkJEe0RNWuwTYJAM+rk0C
02BTZNQRSmMqfrJ2G6AbjY4PRT3O758E0eiqAn8LqX+Ev8lUprrwWhXppzbl6De5
Scko+22L6qkoXlc6K91c9amprJhWMles5WGD2ZAKwOLwOU7Tsaf6pDnonl9WrSUX
Q6qgiRp/FeF13reMaW63888gFMRqoC1GX2mAXVZRGjsxrg6LlZVs01lC70SaGrvb
Qfbp0BCNfNc3HMt9QZKVohNLHL+qhS26O1+9m3idS5Ijb+xjvdFvtc2fZSOYzvpx
aH2jdsrMkx5foshKGCXK7CuPDE9FTlBjHrNKX6mZamsDJvrqMVn32hoISoG2QYfJ
PZXYKhm/3cjRsT9jJAIM3y7bXrenaYNBog91GxcF/V3F2kOT5Q8BHqVYAvH2/uFK
kTBUinTkAfRfttQbkkLOtT8I8fiUZ/9UHKhq57Qao3hVDnCG/uywIWTgKvy+/TOM
P1jnGYMTmaTgogzaGaZygZuEJqmpaJPsLgsBTDQ92vkZ21G6hmIvF/H64WnTwwpp
B9wYKOniP80E7jJ/X1iGkjOBOYoVJdkaaoQ5zod2X1OqyipRaB86CGpMFFHi40nu
wMJA0z53oC9rva2okqc8/UK6ykc3ZOxHX/I2VyTnJD2IsZfbnXaWYV2H1zc/O3si
ZmWywkue1BLWq/fkVHqZUyMv66xQml5+2wtQIbRHp9I0U7KqU/VuzfQ0ULmi5V8u
o7AWt5qr68xpmlfhTYTNDCm74/JcKs2F5+yfi7+xZAl/6qGKFJE8v5nqz8uafeZa
oxi2cJVBua8PB76vVUr1auAojlGSwPUKSwKpJ8t6Gwt3lOSWspcKMuQMruQngynt
cNl4WJZGIJCCrXEfoZJSLpzH9/lzsfBzXEtWycWoUhi5Q0Ipgm1WE9WKlkkAQ9dS
ra2V40gYVTdhZMfp5BXt2eWs4LpJCRcLMhCuai8nJTLEabAZo8q8NnGvDo3BCMDx
NhxtuwzhV2/9Z9QAS5zkjEo28P547F0Y+2Ov4jrQF0SaKfpFAh7x2ISEqtLdA32v
5fmL+WiHP/U9ufnS2Y8bB8KT/3seaPZFQi3RbQDd3ItL5fCmi7p+93M+pcoBD26E
XyPRJ2iFyXtUn11RxrzBx9f6s+Dwy2Gf1r464h0Y2YW61NdDkl+p1Cc8bOkD5OPb
dRZqjxYpuzCk+tCJxk+LXrcmU8Tc9rdMOMg4/iQsbjnZHeZj5aZ66cwlKCxbzsHt
B+9P9E0zUtDXDUjK4Q1aVDbWbB5dvTJ03wmjuaV4/efwTy9HCrSW+5PlTUEgMcvA
UmrwsBMzH6yEbCQt3q3TE67bcHkWwNlQhxflKarSw+Lr0syXtguSrLoh+HXq+fij
CrDaogRJJevHNmQQuDEL6w/ZR/CupdCXZAh66SUth4qifyqE7Z0Ugoyv8Pj/JGwh
E0EnaUsfZTpCkQSxkEwiviWpJooRnxdLQBOG9+BaikkvWwRjqNI+Vlz7rq+3HeaY
//ishue7DGGnWwaSKqoOTPY3PIWePyFeGf3o9lXc3iA/pTeJzSuNUTWZsfApVZFX
aT1vWPATtED6EBDxgeW18HUJZo9AiYjOPWpMxcYBb3JcGYYpcTLAomBWBNaiSOX7
ERP37UHuaYVGoNoc4R2aacC00G1EzHVVY9OMuvIQHmoBldO/YVeX4okKJww/xWUT
C96tsVG+iBK+iPDk3MBUSeMhbra2rIamENSsoh0GFrgSzva6dHzWZF+z+aV2adSE
LASufrV0vUXtVkMycvurKdOaWtVVFUxnXzP4spvQx7XHgM64W6ilAF74VLZ5Atp4
lUFmGDz+6B3urhQGEgKg3JiRUsLl18C6nvkoyBaeHVlQreirR2e0Mscks7bzzTw6
ITLpAQHKTR+HQ5FxKE6VLAJviV1gNO5c0SW1bcXkqLCXN2z2uXQwYu3mzwgbWKuR
m9UrBsI23WaOrlKVNTr1ncayz811tFfzQt+h/aZnkTnTuByfVIuYxT2gNgExtdco
TbAXTkAMaNO+SXlOOaxHMLzO/YOCSqABBz5Vn35nW4ocL03+t6bVqTUR6WY7Mtma
Wah0VSLMpNw/Uc7FZ0eh4zo3HoReFaKWqagx6HIFoiG4bRURjO9xepwqTREisFoQ
2zp8ml/I5hUfh8BaUHBkw0DTpufT2IIwXaWsS3t0GmA7NE7l4mu0tTKXXizY/SzE
8ffo4/v5G44OsulTtC3Pa27DgWXv+8R2cm+j6K3b6bPVKMl15FB0Idk5vBn6TgCw
VizEg01dtLZLKX+wewu1C6L3ZMC3kgWjlptqMilAvQVgeXXg6pfH3KKEsVsgY1E3
up0gjO49lBeYaranK3suXgWgFVTd3cj/cWyMvM+Q6ytYja3LG0+JDo7ukFGbu34L
jyLG9NDzejedGMIMGePfDafBw5La3+vCa8BZMPnLyJSC/BT4k8EQTpzNxGOREgLM
nSfP0DcgLgyThPhujqq4TSqlz35SKPeGzMYxNDNnORZXOX7pEi3qPpcCALnJPkOF
YlNW8yMMIAAWJii1hw9PAR4bxJ+Jg8fmUDAeoVozsuMd2G77WqRvTILmHEFV3Yov
xgfb52gELsMku8y5prFBvQWs9eXQ3Z4qwboVWTGcVEkQmDKGNbsFB+ey+NS2AwDv
K5F/bzmbue48G8teITvjELzij+XNr/23bBvfJp2P+zWv0BS40h6cE/+U6VbUZqlp
itGQU3gZ7fcBBSplm/i25rwEBaB4qc4fhocVFJvYynShxjyQwloahos80e5ALQj6
CywFxdx18gFNGX6jAqKe7Y0sgacrQGSbPR6fTj0QucQZyT4FiSJqZf23cmxm+FSQ
Bz0urcZiIgtm8P1SFsKyYuuTbXnQlzYuRhk1TL0+tBt48Pn653t1BYL8gKhMBCLL
vCBQ7Elo4zyy2B+FvpUtjspvoKW8apmU0UIzfZF9IaNjmL3WRtlsqnga+tVhuObG
SllWl2BlvYcshLvEuNi9lHPfyDUiRv/yTBOlOHUL4ttkvUmJtR6oFqXXwmAugOui
pu1A98H4sdJrAajIxFz0E3SH72I1z3SPCKGo5gh+4Jy44zwIyQDvaz8EKclT12G5
syv4CjJnjK0xangBJcLbZjPFwbOpZmF7yeb8VCdaeFJVZ6H0AvfjTCcdc7V4kY83
S4EvBYnjo1EGFeo/Tjyvnvc0fXPTiK55F/LbvxtJ6mr4UeMRRF5SB9khzTPsy4WN
KGG+ebsnvf//rsPc9fgLZ9PHWROEIbAlylgSqQV+ZWwFiHL6u0nUgpmV2Mr6cPFo
x9k1lHLmNAiXNsi1GJ+l5nhJ0zPYhVDDsltfhh6x1ViESZijot7en2414sghmlz2
BKIbWuDeOtEBpQrziruoxSlje1x21yPuvaH0fRC/zJ3M2so8K2sTxxYLkLu4VqTQ
8pE6L0LiVb0NavrlCONUwY8Tlq+x09dqM/LSadjHKoKkfKXtWzwvrte5AW2DXR+k
JgvStOdFCcrK9hedrlO4rxFVLnU1wra/XY/6RPZyhWuM1m7Gus+G6x9cJWYtVviw
6UW2kLZ3c8bfKdbNq7IFmV61fNbr7ngSMaDik29SjCRPd/7ypkS8vgLDpstSjCy0
zcP2KxbF4Vsx90Ejw/NvnnbpW3oiGhnu9mjmyxQwBJ6ktZTCJwgJRBYt6FPoKw8s
ObOwQ3esvCq+IXQaSH+rgGewKRgL8t11T3jx4/BStaQNyTa/twXXm/Vtn+BRuBVV
Lz4MZDUo8hssjlvtGsiwBM+22eoVizhZWRXUQ4xLmBkPWY3IzHyzRREx0xV0pEqq
jjcmzpJZyfu5KZiiVZuWoClaV1DNFr6OgdKzmrrW8v6RWC2S9QRc/dJxDsYDr1y3
UQTOUAq58Z2v42e4yJylovs+XlXtso+9r7zQ9ydZG/JxORUD5BzBLwRdZSc+NVDt
zX6WJOTasfQmbSH1g6qfQm1wLghqeKMRIjKHTkU/FMDnM2UBzKQNiaXJc4xXLCCm
ArT68QzKiS8w2jVu/ZlTwd5EAu2TIx3xCuG7N8T8wLFutili0obryFkrG3hSv5rP
ELDwP+0ZrGuDZtfHEvatZauVWbYesuKoCP/5TLKCumFlxXJuwUoLNbJUVLEjJF5q
5hg8A/O22DVg9EK8sXVIVP7rqVFPEgsoUYHaxWXKNiqpmv9JKllT30tludMrWrw/
1brRDMVTLJ/dNXrIKKYKO0oX2qGLpr6LekZ//WO47suX2RiyeRG5jwDUMCbO+oLy
9wkx7SMsfNSM0q8PsOpcZQmwUXvXg1Cib7qNyEGm9P4CibcvNqKv1WN++q3UKK2b
AcKzS+KYgfuPW/G2cjFMeYhjQZAfEEBNPhq5kkchVdyJR/y3cZFHqJp1aJSkht3H
2kWU9qlHQahTLM/JTp1xi2z+AwUUD6BvShbrwvAF4m7YDuDALzmFWO3FFAOVtY/P
wcl2HsYeDcfMF1brpBbtNnwqt68GB3aHSCh7bThhlo8DdEewaEWHARbNOV09Y3aQ
3fM76kaWi5kQcbvD10m9f1yq2gqZjPzFHV6ql/FiMkdC8K6iUONbsNUA4Ra+R6Tl
Rqoqw8Gmtw6p0Ufo4lm1BlLf/CvQg2BM5l/JEoCmAPO576YkFhpO4f16q+bMfiHw
ZvkSogpthT8GS1MYkzGHgfWVv0vHYmrSHsS+9UnIlEg6OSr5/Mbb9X5GXj+4zMgm
f1EwB5Po0wsWbavDvDTRyabPF2BxCxTACu3WNvUqckBVTUtNsrocptP2TLD7lcN9
R9AIjGVWLaV7zfci0ewJegQuiH+x6nFqumOJKJvxXU1kNactRMxwVgPmXeWZPJMR
BJG2iHfMV9x/hG9HmnGkQEtsAw1g98jEw9i0ua9EeQCfEkOsQbUYDJl5kAqNUjrZ
A7YHkp/mJegal/kTBJ82JTQ0C0/CkUF3JuAfFa2EKJIgl250ftAhbw9ZZAnC5z/Q
XnnvKgW2OMweSIbjpdIZZBt+yVfTBdysDTDezY3BneuU7Vew6UScC+HfDkjzpg5a
HuRRJMH+rVD3a6W8U1hUhx+Dr3i96onSdJ0B2/j3C46SvTleblWc+5R7qtS8QYDw
sEevGsxZfuRPAwY9Fm37IuK6msWtbwpXZKfEUN5TUEnj4TN9SV7Cm85HxWoDLOxW
QzULcPyCQ7XFyv7xa/5+pqwa8qihKv4Vu8TBjLiLK2iFERT9NSCn56BfKymdfyC9
QZSgwFvJ3wFMLLiYfvMvIlqCKNSwcLXljtxIU6hBXfD4o0QSckFzAYUiiPBTMG/7
8gbe+d74TQ8bc3tziba46kmtvH+kaiJOxnJKy7k0eDJ8WwM4iGpyMUAytDdqudEg
d47La5jX8iuiZAPxDnXAB4GyDD2VFqro9o5VOTjoT1dotEGODGuFGzn/SOlY2/y/
83KkAh4S1KD1edfiTKeexxNZxwnplVpjdQmcS39aZB1rOSuNMDqHMAy0wJrn3oDh
/I5Dl1BWa4BT2gcQfwj2O1FluyH8zzkaw5xspttHsa1gb1Qp5+d36b5QD5oVk9Im
N4HEVobzPQleH17swR4iQp5lZWho14oqKM/QCLQqhaYWxRcCmbpJwqCmKyMytDk0
1+CXTH4Yjx3MvDMvZD1TD/DpJcZ6FeMQTlNo0+Pp4mmLzjTSnJT35pp+tpXELD90
330WAhVaiBqDBdVFd19y4V7C0KCeQ4U8vTbiyDuzqM+o/AcGS5HOljIREiFviO1S
VCyUAqoqxs7sjOSKgVTp0ONOUcpeRjhC+/kROmAFe1GXI3Bnt6kzbv4iuNdb2kjc
l1Yo5vqKfHXkER9mAflNntCjqBRwBV8Ui3NBZNR388j6UQk2rIvZmybZFwYXQ1o/
Zz6VV8yQEC3SWz9sj89B00pvW936/pvma67DoDLe4REXC5puTlQ0+xJ1vQ4PVekI
cd9ZsA15yO8fs933bdvkxsakbEApzlO1P6/JB/gdkqLRVj199puVfrHkpr7iOOEu
Ee12SmEwHs3uVeUmTScBEI2eSjsmRXvjhVQ4Jqg3h804R/WHv1O26w4wYdHN0O91
S59anwFI5x/bLEV01LPFoVepbkEXC8pixEDmd9vNRMUHPU4Jlsv2eWB/koYNdKge
Cqmnw+YwxthnvFg7zPb03Sawed7aamsx+ubKIzDZroiy+6T0bSDrzut/jpOVg8AG
19tlDfTzEtJrfT9lEnbaBH8WncI6qet13qFX8M867UIquoJXtEi+SJd0nm8xyNl1
VRwjV4ILDM2BGc+f8g8a+q4qEVjY03SdW+F7/ubEZd/jaQwIoioGZqOkqrpxhyL0
g6xgOI5NAN3L3lVRlUCewOn+BGirRGuieJm7/0OoaaLLST+5UcHvkW9W0Obar+s4
9eNu1lDoY5mVBcEwHCVCVK+IbQ3nAC0Q6iQwUC0JRHxUWFwi65VpbTpxyLMNMO4r
1ZffOqUJW4JVKevzM5I/7yyVof1GbCqHBBbSs/FLKkR1muHIHYafbpafjCbFqEf2
mVdZ1XVrVZalG8xwo0D2dmvPpskTtyBZG6rEtDdGWhdmpe61QIyIPFEl63pWnTC5
WzgqwXPPeKSikuWp38KDTmcyVcmTyOUHOuPCN4Psbb9MtkBa3jsevdHMUId+TNxI
vMwcWhjzBQMiqpri+BOJdTZCPudwTfTr360GFPmcJlDfeiAqq7RBNZYtCoEa4ZsM
wvqM7rHPZNsprJ5CH5z9Hnd8EuS623jKDojY6Z1go54EZP9wRL1Ffzjm0VXRuKdv
qQpP9I2CcKVH4nhM9wQrwDezf9c8U6axwv4MZsC5IJ7bHyeuhtrg7rZVIKsomxUb
/YCU3t7hGa2chdaQtq7gSU7laQGz4+6dGLoY3id2JqZ9g7PVxNeYmSpC9hzkZ6yp
x3YAli8Zs3QDNei/evhil5xEkpONtvBS3JmFYaMyLBi7GphvJGb/iCUE4JkYwmbd
lrsWh8XV3mNx+sRO8hFNfbC5I4x5VNjwaG37YOv+Tjla1ePpnHpnDwzSOYSUI406
A9O2wMGj2y+JTa0krbIRhEyW5hs/1Vw+6CfB9KfT0EI4CkLtYtClZxhjLrfTn4Wg
r+qaCXdTsgUh7YBqhy9vkbIFCTW+NKDgLS7T6Uql/a9ji2ZPhaBppFB6gkcd3IyC
HLNKvi7y2nWVOafEbb9+UgCbpsxhjXA0TECgviSgCMNJ2eVoxyGhWU/NiYxqnMZv
e4WG6ZtKPgo44uxUQDVJlpG2qZnZjPrWgooWLnvoIy8eFB7AnMurwmMke6hCZPTE
Zx6F0CeHzuD3atOwbecJZUbzUZWMm5+AbnA+vzWUcGplGR8jYnrY5UrBFlhgix0H
89xfmFRr3njaC9vfEiwbxhVR8GSulgm9t8XndTaFPZSItZX4xnPTLV2QawoIRjST
lGca7bbUtLjOgF9+Ll5GMkUDXfXaoPExCioV/6E1njixjRsY7vYYlZm2tro0uED8
2ttIdhsjVcqmw+yJZB6DycbI2BuRwy3HHob7TCYxZW2zJ6QnauwSq2Iu/tgb9Y70
mLGdtaVDRTriIWYbkkmHJC/DQx0mNskg/oHByTKxumREiVJWrJkp5pXGWghzw/GF
xkBzVhEIBo1iFaWicFXR60gInTqvyvTlQBhNIlSh57LnrR3OW3NEEqoYXdt18uqC
nijmtzrRiIPZ+W8MHFje8jV5syJZ6LwJyYiWiBrMVZSzBGFcmtXW+g6f/PyO9hFf
+Siz5+XOTHe4XgyUbPF6nijZ2eu44iOGaOhLNf9c6H+z8Klji+RfPb5r+TAJIfNc
6LMxzx3RvEwCb8DKZaVYXzaxcZsgDQnk82VyhBtJJnKOODnauK1g5iOp6qcOU3hf
xmCE/P3Ah2IsKor4eXahFJqMwOL5yiAZAw7z4UMOd+hMRng95pPObSz2TvbbYFkz
J+upAqYf6iEKsdvYStypq5tnnsKSdi3vI+iN5Ey1Z3SLUw3f1ePUXDXQXJ6NZYl3
IijfmGkes8A3SzHdUgHVTA9mXHyBizIc7GXj8K4YOcK5GrOMLhrZrHLciemGVOoE
a64MejvLr8tKRpMh2fTul6/TkpQ7df1LhqWlpTbsSWeMJoNytbRjDPH5p7OfF/1w
VOO1rSio8erwKNDWsGkFi+tRfNeTWDeXsc04rC9N6ydGxEUrY3zmhnfMidwjm5by
J5it+SUjB6RZWrrF3gP7Jzabv61D0bcSIwM0ZuiUKPlu4NpDlXC33F454ktOKu0L
uHoNw944CGNw4uzx5YhNQlI+Bn4JveeijUc6hU9hapRa9RVCeRWeFf6ulWMkInie
OUq60NDiqJszVEn2pKgPkvIciVeXR86evGd5l4DR92p+uyvp587qbBxwb0fDb/Qn
ycGdVG6loC5toGLcIP9z13+9plPYdEkyehnsvIKQxg6jaOhij57AqitDCnWZcEul
pqk2/XyvYzdCHpKwVVdAcvT9ODigkV5k44G9ce3tObnMtuvzsNEPLHxBtmke7tyo
UIJ1hra6dc8tGoIc4i05AMpZlKage7/NQvdYe9RmMcd0TVPcao6nLe1w5Wj4DGc5
aYqhY3fGI4hTjB+W7U/YaCZC4HA5fg48rMX9Yb9nObLjyg+DKwK/VBkEC8jbIQa8
AezAAFAYsqfEw/lCycTFSv324AE1IbmEA2+9OiBfvmrcWkPMLPehSwBloDDJ2++5
s2nzVueR5RtFOE5u2sgt9NVVBZBdmSvKikBfjKEDPG0igp2Q+TpVdfIlUi6Cda5E
CnjHlaybdig5lw1Ct1qfnlj333XyQHnX7inrGuiP8b+bTvsOY5KRjy0M+bL1Vrp8
xm33CXSOrOi3HLZIFnY2wg9CMON+AqQ0dY5pv1m93gQRzgoU2dBMyYBE6B7UE6uk
CbehjRYLkrcOytamLo8RBYJVTL4hfr/mRKuFCaSjfKG2FamQ6SO8dtZ20ad1KslZ
z7qx1q17iLt/vnGy7IOCskmV04TptyFvHuy5wBbo6wX664bEnUQwkB/tYWzwVqW9
ZaooG2bpo6TnaZFjQuUYHpBzMMM1sN9x1mVS7/c0Yw0+fIGxztpeuSvXnoiuc8M5
B4fj/qmMSL00BxDYlPcz+zriWWMlu9ZYMg2gePvIvz9OSavBeUu7UPzBzeKDF7BN
YNliHoeMbA/hGDAxwA72TasfzED/EJNBH4rIla3QKmsrsWl1bPnoP+yf34wMQCkJ
bufzYWUJ5nbrYhTvehRJUHM8zbE4MlqXFXJU1QrtTeK98Ur8GFcN3gA48kKle7eL
KYXi8Gg6Ko95uUzxt8k6TtB9tAUTLmKdzJ1jRh7NHpYyx22f6Gl2m2fvmEqkXbuc
U4FREUIE+yeT2romNlup8wgvgTI+NAomdhOv9MiZWl4ZB1u2ajARWezF7U722qYP
QpLzuw7+PLD3DeYpoOaUXuO6Xc6S9grlZa3whAdSUVgUyl7n0nOL230zqXUfZcwu
uIW44k90l4NLfbuN75agtOEY9BcQzgeJR5OBoVsfuDQMXKpZV9x1L5DSypf5JMgt
dSlw6uGSPS95qL2YGhsB7YQ+Py61kcZ3ehmTHLxVTWMsycCYZT19z2MlQJcYjI/F
geM2ds+aGAZhOTO8GwMtOidqZYp/5M2QkJaP8XwKxpaH5gZfPKuT4jxIaWrzYNQE
BnRETk0XB64mGlXb2OpkKYJsOThW6yzas9EmhLGLdLGt+I3eIkUQl57zynr2pifs
k3r1Pnzu3SjUNv6ZWXU1KWr6il8DwL3n+kTc0JvoUwA0ZBu+tOz61O1xYoYwp1Vq
7l+LMpf7HCV7ptMAm8CtL/YUPHgQkaoGUnPlFolJhwjAOcFihwCJOnrUIZbPnsuU
3PHBJDtBjNI6BQVYx9HiwdQ56iwhegAh7h2o+JdVtrxoglrZyYUPz1U6QKgmly2r
inpiZOg+DFFLdkaYjcnMg6XKu9p992EVSYBPhgoOHmDILW2/hVB+QeUOQ6Pywml/
ZRI3V39MljaLbHd4vhZ8Zkc1I5APztWymGRKdh6IjUsVAR6+bydrZmX8CkDCxr+s
ezIcwJXFy29LMsDNDrQo9mJCS6HueqvRtHz5cmy4Z423NeMXZhOtqNppvxhPqVfY
GIrsNJqjxrQW7Eyx8kykzwELVMEXPrR3Q8PGf+f1Qd2fI/gU8YDKyPtbP8jzM6i/
R2mBJsn9DcHHkw/k3L1bSsosggn/RkbxJqbnEeHFZE0QvK+Z7KMvQQzwLTvhRCyp
cJjx2PgEalGuhsyuGOff04NCci87LPiV0UxBoRnC7Wq0W2/wGu9zWh81ygMab9r/
NL81Q3qaqUMvaAmAo4zaY/maor79bq9gOHpIjGMmss6awSYk55U96THMcy1qYGp0
hCmkikrnepGhFnhhwiPeGXsrHu8kOufhezOWK076qdVaQS5HfsZnijKOgve7YhCi
UzjDl1iz1xbY0RBKwLlK+WkrCzUf0B01O7nAHlCKDcZLBbqkYSK7T+lwT5AxWdLs
TUztfna8nM//HaCI1JpzFgjNkUM6/zQWZ8ehHqgsilfn3tOxnZu+HPuXewBbrNvi
AL9Lkphg8SKZnp6bpVSTkLc7CO6TkpE1YZHHufWFpKDMeJbS7UBGeAC3vM2brGml
yT8MhF9+oZqQPsI00Wc2QMTjIr9Z7D6gDNPWPDXe/714hk5bs57H9wtrhaN04Mpe
JU6sz4ftVTzI0NuwXzv+/d5dWDcYahgTP/u2hKTHQ7fBiaUkbIqwr+wIiZNC+KQv
QHvU2ADeLQlNnBHn6qqU4l46+obESnByGXtMKsr8HCn3jd/qmPN98mHVvLN4bXc0
Hw0rFh51tPYTxehwzN1rgk3B9A+j9eYQctQWVSzfxNGOBvOcHTEND3f8fJ2h2BhM
EtTAj0zcGMiVBgntrUnT8bgrLpYVIgJXQlxv/LGCSBjDle/vDLTzoX2MZL8LmTXl
2Nlz9J12tyoLNmYDy3FQoiiNEACkDsK2DahkqvIOJ7dK7Hti1Zy3xZ7i3qSnogt5
kPCbPE2YTqgMBhQZSh4Kq/DnRQ+9gqAsOU08k7zw+f7TZzNybtK+ux8PKlr5SoZd
AWNCKS5LZkoxR62w+4/9S9MIf65civnMGF9/TX6NZz1sRKymzeasCnPAX5/DdVaS
HhkByvw4U6RJ1l+ZuTDoPoOICw3wf1ViglhDs3UG0x+sae/0FJBDPC2SGq2VWQ6X
Eug03hE0oezSC4tIyd0ku2H6L1ocbpJuYqAXoYD33UZzRSRWrpauctp+RGHO+mUT
z7pL0+h4KQqRltOBQUWGt269iICtJdtDtalDL8hmwZyHjA22UUBssi9jVhPR+Jvx
I8fJ32/N5/joRzp2lgyo5IBngeonbf9SN7qDp04yiM9e2av5fCnbosMZALC+bYxf
vKFnZeslEH2GamO5vyecGxGJr9zxKiT+R++oQcj3d0WYgrLVGX+Y/xpTbgFp2qBq
v9goUdlXa+QoxlKZfBbmXIy1Jg4BP9Eifu0vXI3oRE4DKy+E/0J8TVbyEMuVFE87
ZwzxgvKGtGliE0mu6QWlGtWvaRs2/gKdjDVkL0gkYH0E2eDOzhjxcLXaYS9m8Gys
P4IzbcI4Iz6P5u5v14UNHkkejS7Ofty717kAusYV2Fzgvwkq4jp4TrOQkwuhUYJq
Pkgt19b6YipdCBF1XV95cSrWew42YXAbhrBc8mUt04NRR8WrGEnvzfPZEGen+suv
SCXyIFhfCc9KNxLLREa41kExqiUOHrCzFJfGgrcy1/S8HfKFCEORpwiIlYJDrgXD
/PPp7eyleO8FKBzsa8dtNHUse2SOfxEW/v21po4p65NQSydTQc+PwbxTto+mFUNF
9KMP2vbJqDaFGmvTIBWOqS7+4LbBcgjZLqsI9bcxnlksN2s/kD1rCHbgOy28QUeo
nmur7XtB+m1V4rg1/zBI1JfrLlpxFI3YhZ9x0g2PPV5FArSSInlsvxxdg7oLOjCL
YeEDyKqb4uohIkrW26W/VNF8xXSHrbYfiksOASv7U9LoDf82FTSpzUQPq7cJMoH+
HROMQQBdo0L8Vn5LLq6za9WKILyi5Ejf/4xx4/yxkK2EvRDQr+keJK9SmrTRq6rJ
9ZWSodLOqhT7C3XFgD2qGXcYCUbGbXev9ioZjU4ij2wfYth0XVjMpCMe8Fkoy+HP
1EftZoWWE5aELt9iFH0Ta8z5pIA+Svl9P1Pkq8MEmV3BzkG9obUSv/TB/y9oZM4e
5L0EUm8VUH2z2f1arn6ENvA0kOBGs40rZ4L+ffEna3T5DqTia0XXQ9NxBh4Z/O2M
9ras+CBrHhw2J6861OyjzQBXD24dEi3enClYtpGF8bNu042C4ytksQLVTybhOtpy
Z+rsDo71KcIgAdXS04KcNXt1kGs2gfjwNoTKgzXX+SnXccC5d4Eu879oI6PyvZQ8
NnUUtOrIyj62VkxDFlRM2Ml5Ib1uIYIFycJs4aXnnDOKcGG04YLMsqwkSb6NsqBh
7dM6BL5M2AaMsEDOf8MoULpGg0WsgyosoFEebzgYMZAAcAfB8AvBPG/ciW10+NLR
r4SKR83QIeVOckS7xAW9NgIktFhDJoT43TQHDOMOAOxP58uFeV2lNpJApr6y0aFB
/O4ZfkJcCEAUurgSqGwKTx/HlNiU8HkIPqe3PQLjUaEbr6UiEqTjTrmfdxPWHPLa
UB3C+4FRa0l6zsCeqbimnclmcygEZlkRkLAFNoRdseSO0zL9GNMvkhaknlrKpcQw
sryil+z37ly6wBNu1rDCeqc66tU5AfDhFWmbD/h/9/Ib9l9k5z+gNztS852vfyIX
rj2KrxfJZFXHPeA9cl+C7EtihRXtpE37K1Qx+3NU1AZV0Ja3N3W5tLgvX+Hxy0Sf
KvVKJGSmqe7YPmUHSpN1Jg158cyGJE4JhH17ouEOlUlfmCVwG0nyMvFnHd1ZGoGm
q5c9YZRGIjSjnH6HeX925GICCXr54FQhXeFXyJ/J5u1Tvvxm6LNHZwj2TJmQ1ZKL
3KcIUIT6YJIgLHd5QflA8/+I2tLwj5BaMJQ7iIPFd84zajSW9bf5M6Xt3/TaK3IA
sAmoUkhfk6ojasqy9KvYoPBld7KN3/uKaPloDNhtFWt1eBSDJCE4UanzlqxMOdAV
WWkkqPy1IqiJM7PaY2bpU2KivMjx7WPslWitZf94IH2mMU+9dsj/uHlDYJRujemn
mxCoEk3vXr301dKSz9yMVHxhtwIV+ZEfFFiN8UWkVA1iIoqRQ0cO04eKSc90oSIW
P0P0O/ftVUhcccqGRH1lZ9T0JV0ADNFxTwtPzUH68t/9plNO5EcZ0hrljIiPrgkn
1LetCiwZrWQZahGEE5mdyXfonEADKQSgx3jQLEbX0RzIeMGGqgBPQ7FHY1iCxg09
mAvolyd6mxD58ucAi7HsG2d4VeKpqj6bmYmlg484LJIUji8kt1UdhzZr92vaYC3l
WbSxj0YWyFAWV/yul8w+0WWo8yVuRxNe2j0HJMe7ZEpUQcog7uFtQ8n6EAusmQbk
qeDVg+w1YJsJZrltwmQb+5ccEsGuUee4FzlXsYSW95EiuQArQLs4cXd3Spv4fDqt
ZO8UvTGrd2xecBf4ObjxPbrscXyCubof6B7AoPqjidm0HcZJrASuRQ0LbWDuVoN0
SDF2wfBIRNnWFoARulTxisIzYjCGm4hXVQFDp5Tv+Y/liSeeG97WjiXi8IYogMKN
4WAopr+Db8bjcOaCk1sKEHqISStQuNomSVYOeWRhtFXfAdbTU7DNMMpaPnZFRcVX
sKBzTVKZo6NHlubE5OkQVI6CYjQsf0yA1/Ha+RhhkruKcTaTOVXKB2by++wT23mF
d5LYQDlhOQHyoxxJ9wOfijHc67+WXUZUGwLJ0z+aFhODbGe3kaJKyTSddp7Fljcn
4u28PbJWVHnEVve2U+0I+GVb1t8ozcXDERaX9BcbKWFgJZjDV0Z/2HuXpyo6Zh1E
UAYCgt2wkHQY3+47hM+BYv0Sz7RC6LHd0atIKYpx28LPP4NeWcG2zx2AwgNwb/la
06cbSkQaprV687wxLonpM2YEEQ3LCQB/2GfQg/LHuwQ5eS4qkt2W36ZsABcgBo9g
hFGpuhDDVcgs5cJgTFsK7jX6bm6p/69aYsxyHw6jnC018EGZ19HPEdKxyWNV0QrK
JoI7Ep4JAkLcFLQruJDFbBdDj73Txn0DRa7QCekdYMkesNpAQs2vl0KN6t32+taL
ISdzFBrCZ7BgesA91SnxvDsXtuyF95EuRJmtdIVbgSfIj0VMr1Rx6VDcCW2frF6m
SAnzNOg1uNnNrPu1vza29vNq5x2/Y2MC7TBz14y3A4caFFHObaQ1L016Ss4sWAWT
3WtcJomb4bUKYySK7lDi4mwdCPP1Z7t+dTIRY1a+yY0/Hb64c3kdJpqF6uuz5foo
Tsrzm97Ypzrhj/Wk6TlWhO+lgKNHr59XK/ppFbgabsTGzEPN57zZ5qOOrogVRPpP
Hu9esIvwWgb0lUXJ+Pa24DqGO+TYKZSdCTgpavmz7HeOvN3ma1miT3jwCDeyVvUU
lrkFeWU4twIWPLwO1PhyRMGFBIwPj0uuEenX372c00aPCBbzNXlXXnX0rfFtVkRJ
+ivMfyvQY58E58niUJ0GxUmMeS8WM08IHwMSucaIezIWCWUtaJyZ1JqmZw2w3C2j
mVOxGQGQZlkCVQeTRZ5nsvCxfCR1vOGGE2OuM8YrXN6ZabGlEQL4gcCYalUDXjM6
tEAvX1vOmyh5KHAsBgXXKbqr4k3Hm9Ng+hdo/YGF/zEjPwRkl5qVXRxBcIC11rsW
/yqyj4j6QlwYkuP6mQVS5KPZmpCTEm7AMIwf60vEpNI7oUxdzFRrXoTL1rkKKJwT
ewB61tRId8PR0P4z3hduCRJVrljagVgNx6LXEZ/Fbl2obD+xJNOOT7GhnXUq5DrJ
CNXlV3r9RlpNTYYRR4F8VTEEbAD+Uy782z5F2lJWWdSfuxJmEXQ1Lj3yKW18KLTr
t0DY15Ayb+XRZnzcREicL1ec93WC6rNZKDHywYivu5UkBlj0mRaav9yzfVfbNlc1
UM27vHNz31agKRocbwvOr5yocNjb3DAHvvW0ccyExitI1LDYe+y76Hgqqu+yVOyv
ggTBmryoPIf0H7+qohrLB6SlklaMjJr13gczKaMGEUg3VzezZHq0tWJ5iS0bXxR5
Rorg08dhxQaxzyxUi007yUDkaq963kxH+zS4orXSyHTSpnCh2LXitnQz3YztWuMr
GhZnfY5JqxpN+smcLVFl8X/SUvwrHB0oy29l3BdJQ30iFUsAAwXIW2gdBhFhdRpX
RS0LnXX7HW1nX/1hgM8aeUu90UCArcCi9AkdXe8RRvGTUkHOrUn/bNjFhHLHXsSq
AlOa5joCgrHSsJl1yf5cO7u21lOXYtHinuR4RePgxJFg5gz6eX01AY8takleDcKd
TRIqmwEm3skCvONtRH85kUHIISTczVgi8P9QRA/6Aenw6IHArA1mLRXWwzngErI9
zQ/DFCxTUNIQVRI74yZWMm2C63dSlIaI3NE6J2iAdblHeNqpKZY8TdyO2HLx1ih7
T/lfmHasgv/F8+UtAP3YbFuflUcrDrEospvNHXpPbS98vURsYnP4rd2rbEcu1MY6
RoV+5748pP/Dp2nwHHmjF4aXg+E9CbTZ9kN8LTfrbcH+/KMsaJ/jCq6BQmeo/CNv
Gg5lpSrovQkjSfH6DEyFWAoi0QoQR74IeLdVsHhP2nvwMpJdcwhwbpSp3BPAsiB8
LCebRvmTbp8q+UsaKu4GRWT902h5IDD6HSIW2cugKdI2n55kN6ZeWQAyXN2Njig2
KU1uVku5vai7P8lhUvWuvDv2dXmnTVWJuRmyeoEB5yFsr0qGkn+OX6tc5nDLvzDb
XxzGypTWRcMTcgFlhYMY+2o1+jYvY8jd1BzWyEqN7bWcJWNegzsniGSu/ucYIazn
91OqVFWCaFt704ledJoKEAVFKbafdNX4AgGiJaF4MRlTwX6Q8g26ezcyYjtvqzuM
uaz9AiXugeumCZjisHFQtZ698kRh+pvUj7uP0gi11FcTkhTPHoxvgFftsNmkzUgw
DiefmROjaerJRnzIICRNQA7Pxi4vC4GzaDcczCdoRoXpAMs6/Y7jFQXQMpu8+4De
lL3IymxKp8D+JeXl9ivtk1x8QHykB80rViDnwwN/KlUKiztmOL65dbs4ZxzjrwjG
tWJPRxySpdP4a38z45WFXjK5dRhNHGMy6AnoxKLTRdO0OSbqI3k3twJHwMysOWpv
YC0hmJJDwb7NKNLpKW9a/oqaVIz1y66EYaXGYGJD0c54leH+eGbqlvX8I56Do5lA
AZiPDfKa06/x/8BZqxe65pDlhsWvDfcjHeEmn9vX3EHaHBnB/pc/qAI9i5h8jzGO
CMyieotArZMT38cCZ72b82WdG7j2CRlgQgg1xOp6yDog0qeVLNoRubznYirDYe88
rMJgOizOSkve+QU91tejFwhQXg7KYi2d0pykpWmQfNx6C8s35fNe1//pGr+08p8B
jsca3FMLNJzm4jrwLpL475qidR2WozBbZV8uCjb6+3wjlJvVx39ATiQaCfrstYpk
FIUp3XW7i5h++un1Mk1+NiyK2wbTFWuHGKrziPZdMXOGqB5IkLsWGQHLNPassIZf
1Y5bqxDZk+7vHUq3rETP7WLQtL6h4Am5+YPdTN+zEyenKf39C3Pit8Ggrav8jkPA
4CUDftiCYSgT//d01ia2fgynxSW1jrDQYUyypKPSCrl5tHWWwzTKE8pvH7OTQA97
qqItb7yzqLg88LbjpSpJRDijq9MDtHInB89m07JeklK/xsbTm3naK8UjZfooNXzz
R9uOazcmZJSeWWZUXkXbXol0Dkjr3ixP5vP13fZJFr1HitapkHRflit9Pl/x3NU6
RccouYr0VVhjIytRWa1/92V0p14QVfcIuCtoYFjl5mbK35ZxJXRXHLNvWyJeDgIY
EfWrwQJlTM5s+OrDtH8tByhBSAbWGOBA+TGsB18eWKSG5WrC7931tlGO6/OR6dsp
QLmw1hbnT2T7jPvDgPyUbAigRZWc2VjE6aA0+w7MYkqLrxesTtpnkmSiJgiZPpeR
6oaiIEp1Q2bSmd31B2Iyd0B0k0Wki7nxQB1CZUpMZQWu4qi210FS4sICBY9WMh74
7PnM2PgiO/9Bc4CO67WKm4ag5x9ZLEu//j81qeoTId3V9jRcIBQ0gh5OYMgTZ523
tPlcfBg4VXKfTJBEbCQdPpID8mGu8o4AFa1NSB/UujyXgX52+qmIR3jAkl5CNz5x
kYbR4BH2KDDQId7UCEbl6eZHz7VAlJrh3Gdb/KujnlvT1YmGKtffyX5XsmkVudED
3ynThMDDgCw0pkXKrHusfEhkQDxAymQ2b/qQBjIce5YpMIeuc3x3FoeUL5rA+pXK
UemlokBP2GHMBZSU0X+uEeo/OswqjgweZmC4keEIPmy9bk60POiO58q612P8Sor9
BlVijDq+jT3YhyIyrPYTrxDVoyxTkJ9J1TahYvmJZERbSp44Vjb2Qxcqz7iGaKJu
+tQRj+h+1UxZF13PeszPHMYjJ+htlvQwlDqOZswV28E/UFBDlQ4wvlJbw1B+HaPt
Ze3Sv1l+s50Wqaf7njHy1MtjfB/Q7D/Utjx6MMmNSi3ET7yRFeAzdghNpCg6/Rss
EK8gi2b87MgLUttJPnaMESOlrF34lj6G8I8lLpIhf0MyxyE7AiGhciu86cfzRMZa
KZOKbbb39bltxfYHl8J0xk3uCHwj4vbu+ZoiSigLzV/4DidpWXDWiAdzNSKdcjx6
OXQTO2jhA0luW/C/mLfOOwuTgnHzK3z1FgeEsWzktl5pgQortTwSaOZVHmLai6jA
MuHzx8ZUlWEkLnzdMeCwdPiRcrAwnJDtDldwYV6n9kMudxd3T/itxU2vEOIZf67J
zEN3whALQrrWFreJbkzDA8qCghC7HjQdWxmJ9JNEvpBR3B6ncVP0Qy5OAunlGjpI
WzY7zFk1PmaKbaRuCFNRK69H+qmSEBa+mYT5D8r77AiyvfHq2v2PstqXyR/j7YDE
TV8dlRPQ80gepmKR/mub1blBnJyrHcTzLmM47mFwZypkArHvhzw5RBYDpMzVHlD9
jtAxlQs8pPO/O7kCcLsOUFlpf2pnepzDTiq2TceghoUeNd6dWA7BdsJrDAzUW/v0
2SF/0U4Mpmxo+vaNBdj0pmYKmmpeASluuRrFvNDYUY7bRT/e/1GDa+ngTdWbkf1s
EBK14PKYwq7Fff9bZQOTweqmli7INHLmEuX7DXtfvcVzQ/yrG8x9ZThb39a41rH9
dEs3FETSQHLZKlzjoeVvhwDzmjWs0aydqrktxz5ZQRnW1kIVaHV9v3A9UTDlv70C
h00cFEa769gzd6IN/EAeYgnmA4qt3SJfiuf7m6X7o4CYzxUZEWJsSaXqVLGXFNJG
5TvVC+8Iwz/bqJJFo/5IoFEq5DV715FcQmPmEY2BUmXth2dFyezyncCRjNhJQqZg
gdMAxjDdxeMmGF0N1AOuTL2lMNO1ped78JX9ut0HtlsRwSgOyIXjQpR3MajdEJKE
TCnJapkrO2Lo0Oj9b+8ZRQtPfiguZPxACKFQy8h01R/Punf6I/YgcBxVlNIMVxkv
rJk715qb8frtrthW53iUoWU2Q5gt0N5r0pLHqNPYCKByzXe1FMuz3jkZuH+rkv7p
/Y7scjtWHbfACIybL2XbGcoTQhv1qWlNuIRYhyk1KX5/kWa2TgFO2DwtO3uQjQB8
5cVqs4NlXVpaFeR3Rpp0Fuo00Vq8/MBH+DkWfnG8qF3PHKXcAoprahvjQasrHUZ/
ViRfP4tnKzFfIYqKJcHKxo5xkTgKjMFa3p7chvhsbCDFCVMZpAdN2ztotiNAQe+x
aodhJwcOucsROo7C18TGxiR20SLPW6ebq8APbR6LLqFdjmhxjn9J7a9ffsiRuZRH
zD3JfeWwe6fzVZWv6eBBTjjF1+UGXpQ/7vCCB14kK2bG5wBe4I+JZGk3N8DGbuqg
vGndm8jpj1xRpfat6IGZPerErwTiAH8ISk/PAU6SlZdYk8i6yyMPFBsORUVLVBzg
zHWADEnVPQlFRJnUJo+ccuNk2ESkaqkryAGS2x8SHecdw87Q9vEV/tDb2BYRZsy1
e4mNnNve1eMObbkKhQ5g04YKjFMVdlx8mxv7ZU8t6pZQO2MEwP02XLEzWc7AE2kI
xcBZjDFg2cTC4IU9Dv35/Bh8a6dvQeu0mMYFJyzl7wBN+iBZrk6Rm6rp6KdxX6V4
ADXAeyrMGtp9F4ibfnQtoRAgax0tTSU4mR98hnVKsbK85XpKLXDyFFNL0hSljH9V
BhxB9cbPhQaoxZUyXy5I0wnVXnaGBhLkH0eBWiaYXJcpMxJHRvI8LWdJh/8Sn+/F
PsKJd6Fm8ziOErWwRiIzoLruq9coQaqhepj2Rwfwa3AQuKjIBQljkvmEApTLmCXB
Fwu45VhMD/UCdmGsrCQyT7zyVe2kN76EjUrcwTVUc1KzAMhu4f3XW/eFWOdds30I
9aCoUnpoKiHkNddeFp3BAUaEavqJwbe+vdYgRdsAx5ndoxvs+OZWTSlOMVWbBrtR
cpBT6YqPS2ZOuBc4s2hBFHCupiujunGpj/NF/GGu3PBnd46PR6sYJ3pNKnTvaMs1
+WAd64iCQqdJyx+W1IuwLnjzMI+M6XI0+NgNdYrxY7G/6JE9GXqFpXt8Y17IYHSE
FIRXlVmbusO95pwhPGV9OZo6Tt74SL5CObDrpcjz9O6JMzFTKbl+yWWur4mFC93/
9gWGCrOLemwyrp3k6ONPt9ZGOlj0vDquhd8TN6nb93CXICnl8P/MapVhx0AL9ix1
+sL4NVJ6BLDHUOVLQPN/MJMNUIvXu6VMFzU9U/VpiB6WBnvFsmNGkvT4DynPK92+
UmcoU0NhlEYVNsvSk+8kMYlak7+IgQqO4uSzY7ds3aHnrhW+EiWvwrfOVxaQGqLu
DAyny9jpOooseXimsc76rHT7F8WGAxGBDsMDZVRgvVhMG8MUllqO9fVWSkahmXpI
xipn3RPy8c+8zHm85gu3iLt8CLdk4i8Gl9XobOMi7M+o/+7uYXoAlD6fN1EDX6aP
RuePA3S+lEJdo6cdmZXrySnuwFOb9wVFQg6PSq5MYQuXoo9KTYKA1fTriFtcDuS/
cM1H1iUo5DbkRAScl9I8VUFh2uD9JoXb7cbgXQ6NFNlB9kFCVzlkskRbIND1rptS
l8myG1LvJztx0s3aZ4i4NBbJ4ft5VEcSFmQ34ZxKFOrUXoB8l54BqzMipRkSSWRn
YGtVzOytgOqt9Lihcj0zgPYIYwLV4Es8GGDzmfNcEB+iyHY4XVK0618SJ3UvDi5m
aQlARyNp/KMghouB1FgnU9ICIcDSEqhglT9ahOR81HPH39ll9ZD7yR1kGzJq4n14
3SZ0XcicyNc1XDyO/osXHykswpA2XFOKzADFsBQImzZCjKcod4/oMNt7fCbo6fnb
un6JriXnMgCHceeKXHa86hrTGsPHaphz8TAcuScTYiQtvzG3BFzZy7mVsTaXYnyr
1dFPzbNrTmGTHxYj+nLwAvjtZ9jDuXuixJj7WOmda7O1dRrluMP9+q4eFOX4f0K7
4RtNyR3n2EFPludtZMfwQbHcZPWnSG4wniLkVCxSssu1pzS1PQIgWux40snatrbg
rnIIg77/G6132FCD5NZSaDTMdm9CjyacV4vUJ71Tibldh0IWmtsLTjhqalTyN/3c
R2qpyXMmXFFPCborKNsZmbf4ElQpqKGY0WI0koqAtRIZOnsH71pFBi/DNtcFrlbT
XOCSdPvzQ//CiMcd5fccxz3l+SMmbkU0XVqFIsTNx68RXovuJmH1P9mLqzlT0FCP
qpUbg+6p4ULvkAaphKmMQdHXcFYfAnZjOggmhov2/H8iTm5XOn8Lu55A7Y52G5Ns
h++L6t6MykU1yMv6BkBfe14PTI6YoLrQmkjRXVLaMid4EvoZYP2JrAyDhKKgU3hl
0/lNy4r5oI8l5kpG7xEkApCiCsTbEsG+8vaydo4TtX9p7BH6WqmhNpDJjjYhEc2K
CYvXeWymgmDd7bgAPgPk/vR1bP0WRx+psefsnFUnA4335iOn0ONhRqqJbv1/QtxQ
nAui6NkJnTAp6vvm88xpwwC7z0jeVurH5SvRKIKiYnEhEvm5B4Z5b3Za4187DENU
uvfU6+dpMLBvK0ZDD8Uv5cg/InPJo4e185oGihHjh3pPPQlBmB3gwKMQCtKEcKqn
f/hu50UbjAqJX0DZUwem19n7wAIu7E/IpWNImDqy4QOZdEnlP1o1DDch9hgCtuVm
vu9+bLgxrk8udswsoBaV4JoLgQFBlJKDW4L2yU8eM64E1y+NkLLoOX2j0clbJAEF
AInIWGzhgAWMGiin0laXXfGJzSxHnqeqVe/MFXQnPRJFAbNqZGRBNnf9GhCXFpeP
TSjpaysfTm7T4kFDlmsOiPriHVLTPWYxt91mTAaAyNLD0yMk9K/CZn2h3IAVgwZy
o12ohkLjbO6dq8zx6ef7nJqTCKGgWhblQC8zQn5KMIkFzrIWr83ibEpgFB2n8Ebl
Yk/Zzkv40fbewgqh0o/MRxlvNMdNGIvwCeh+JCj/t2toNRco3oCA2oghDGbq4OYM
ub5sP9zBTl8RLh8F3AyLW91rt2CNqsEfJy60rsY5YfIQz5DmL8elHKBoC3yX2tzh
Zcm6EF1Kim0o/psMdAV/f0o/wFqfcxY+H2TM+vouhY56b1FhJIxA8i7OmKJnKbYP
J6kJFN8ssnxmH2qb+TtqPBJP4G3Ib2ovdogyNMckzShz1DHMk+sVTMX5skjfwbPV
nRqiavuZ0RJ1p0YKHJqI3/UD/vuSDNuT/DTuMukjX1qQXODxFoBd14Iofy6skLMB
wDZXpC3HNaLARjKYNwm/yMWoS7kppZiixgv2IgwPQ/svvCSxBdrjrByUfBUej6sE
w1yBz6Exy6X4wdyK6/xPW/LZrUykMIUeKgiqaJNrJooVR2ks8APTx0vo4PVPFzIg
9PqIrjHJHre81QRUa6Yq74JT0u9ezPi1WBYZU/1KGQpMIFGTTomyj1IUfVBXSv8r
PcB2wsKHgWi8SSQAuGlMf9RXXpr5p0Fa6OvuG5fH6DC4emRrrOBhR9oyJmVPhIlr
mkJqBjv4/0U1C2S5EAQetVbhIN2X3Y+UJyFzCE+P1uK9Uk6SUWs5YcE5UHLHjVT/
UZ+oQIuXgqUxAE3lJ1rftaUDPVcCbN5pqDqSUgxWqco/SbPCluVS8GB02etRKZuL
6SjzfBqPddUaTr7EsYz9ffaKMFZ/3W70fhjbdhjwC0gmVOvEyX269jPs29nk2Gsh
TTDNJCpNxqb8sBgojOEutla03PjugkZty+q2ePS5mGOeGIzHqB58bZMq8PX5hbjs
5jxfcmY2b6ngTtLONvyTrzQCWvZos1l2zm1D4Vz3q+qrIy3VNrhlTGxH6SeVWmMY
H67QaaFDlOysJGkXVY2ha6IRGpfxkkmgRv6b4QOQo8A6swwDcgqMuOG8m2/r3UMf
UIQ78rFm+Z9ybgMMg8Il1dC5R5gxMoEyRqGyTniUxXcLrwngCi45LOsj1D+TsWFM
mhaCnQWBqkMvvzIlUEGJDMrL86pEY1tfRviCzAkFTePQyRfTZ0e8XdTg4NPffe72
uvwytHILRPFD1fiKeOGmHI84nHIPdq3BC4ZOxEZchMwPhVxgwc6MwqLkvOcQ9YVP
fp8DDyaZTJliXI3IkbOzjlc9I6aE/R8UmHaMGpdSyi3qnIXW9oeBdUQumh7PwEbc
HFxcsL/GZ8l9FeKlafQ8cXviQJjsi9uJKyk7XthYGFb5Zo61XVslJyImalAJdoN4
l2fSNpEBus6nHR4jifrNGDowsvpXBllInSRXLy83sJEMWKyzbjeNP0Mz/aGiMz/l
HZaKTNs1tf9eJXrMS5EoG/SnSbh3swLGt2BGXw7KjdsGpBIGjfmiDC0d8jblt4eC
7j9EWdfy2sxJLLl8q/54H38YD/snQxvMu4EYrkpcKN20lrGznFrdXUCTZ34i04ny
r4mRME4zJ6uFAz15J+bikrK6y9Ou+8DHCAuGRFuWl+84jl5xS0MlEcx9GJX8Kg6o
781utms7CY6v8XAMHb1wscmQbb7HIxCLKl6WD7SlVjBNwPDmal9+CyVo3NZxswv9
0eG6Z9GDjv8Ay8OdErg4W91ozaZeF2SeL6QSiI0hl6joOOY4Jm5aAnVlXzRn0XbY
H29Lvhk5XLmR44AlZzhex5JGGGVjUx5JgC5pv8D0JxxeYXOlm4vhq3DjPBEh4MOs
tqLj0OXIMZBaJyiGGpJK+TEMVXzp5aNswFapzFfmo8gDXdqfrf/BUYrv0Nalxf1a
lJSoyvgkE8qNdcS3bSVe7mn9Ju8VUpdP+M9rJacG6u0+vyuAWnMlL0x+Hh73RJny
P6XolrgjsIy/phajNDu/5/EOMFDDCv4OGQHAs0dw37ZaHYBabYH2iMI+FpZ4NttX
qVYpuCJBL34K2qXmVtPqwKumvI43JKze83PMmGdMnCOQi09qDonTD9QRcNW7RWPD
STBIlLzldkQBK0vDYlA0+laVkZgWl4ykwvgPs5fGfql9Y0xX1TylfEQbXmP2DnOa
6YBpKimhg2BiI+Rzb51/Yg7kHRJAKjkkso2wqkhMDogTtqCOcPaK5fVYl8s6p39i
RetS+k5UeHCtAECB/JPvMNTCfJ+19gQE9c3r6J0wPUZstMiBAxpPJBD1HjXuA1OG
OZQJuUG2rRtbnDYCkBlyXsVXt06Xj27RZiDyPlvrq1QAFXhpBp9A6UuUtT897+eU
7a+3uc6L6WwmRfeeKDOtqY8Jf6XOLHtXdoAvBTMRNgxMi+ql8SxxnylZpRozFTMV
XMcUDEXsC2XT455X8x8A1f+Mp0gSce6fWUzCjVD+6sHrhfE72gtz9XYRCwYxyZhQ
YT1cYfrvqs7jfxAVTAd1kPCP7HKRR1uKgMWqihRPiK9/RK+eREZvyww5uC0D5fK/
ztObKCB/LBMbOXAq4vgSvLpqc1UnDy9pXquS+pTpoJW0Ciy2Gdf9yWdqO3HnDMfe
Iiq+hTDZBWVEdEjoWtWml8tV2cjSu5b7Joz+0kwxcRxvfsGk+4z2/pROmi0aAynF
SHKXgdDiuVIkVToD8d6AK3Cr8SIPNbEOMoSgVi0AqKRo/d0HZzGNwitp9Bi8Zo3A
Dtm3iYPBxWZqUjl6QHx+pZ0iLprDDZV/X8reUQegWNzHkwzBlIpluJDZyZuC/x9x
5TyvHdgThREkRmWcTIzS6p4t6+O10bjGob0VeeGNtQ5gpwrPpP+8OGZhX6joQTf/
aIWCKZCS2/laeOqfRfWelX9m/9EVMWNpdG02WuSg3QMlWu9kRjhE8lXoRgvWkN2a
7sBWafDVPBBdb6tEFdfGJ7m6nWzcQu64KGi0Mb7WWjMJvvinA269Dc91Z8IbV0/b
VO4OIOXXP29zLR+LD/HRVjNUDOLO09iPrbEP0VXCetr+DxZXYLsseetE6UppIn8W
ywqycB2jOGyZFFjms7sVXFtlnmQYIn4eeV1kjyk8I9JMog7l6qr8OGqs3Bhn8YE2
R8srd2/iAtt38QEm5C9f0J56oU0Ug6+h2J1AVFMZ8ZfLYbCbcC2Gk1hctuQaDIIq
Hu9JNp2xPvr1OkUlIwaYsHccYvz2Ln/jT1ESFPaQ6afut0PGm9b1ilN672MvpUAF
DyzvCevqaM5uq6PrRyIOIaOIUhbG7EpBblPaMO3Jv06MC22SdEfiG7+zELXBrwH9
081eoexeOF/TRmPHfl9hD/OIZ7bUPUwn7vZ+b++YuyBhDLGS2DKkUCQVuUG1h699
HC0AO3oVrZmX+hjCofwmytcju2GoW36947BwX0URDLEkLHS8i7+K1mxBX97mE+JJ
WEon7EbDpJML+hbj8dqB/NgjRyO0l6TcrGFU693ljq1ZIPs2SvrRC9ka72cWfrAj
Hxyutg0MtJURdFS4yfOXqPHlhijElicC5ZlxV3gBmU/Q7hI6rbjz/Y22goCqAJin
HfZtvthCaiIQzsA5kxWzxRRFkgjlBbPX43z0GSEoOYeoULVFJZlfCD19JrE4P7vk
Txrh+/i3MrQBxQ8PlNnxfjeSU4hEPHbHYBqhwJ+br2fZT33SJCa/futCjAxmEhfK
DXjo1vUyabziud4frJMlgv9JkwdncH14SehacLgHulhL8t4mrtnEurkIFWE/azPI
YM1PYiI5MpdzulcDZKqCCL9nRdmc4f0XMM4X5CLsXGBM/Pu+LFNIPB6/ixbLIxPw
jnfcDi7F6CqtQSF0JcqoZ6oXQigoQdJf8T1GBBwibxw6mnhf3ovxnNWovfpApgJQ
9sMLpxLlu5vnFkbIP/k2VTPBC3Vew+qRMr/u40a2Ox6I4cIrM+OddSJAxQEWUcmT
GwGcia08NOKFpR6Qrxx0X+gsQCdAWePK9jqUPKXl8BeTm7gtiqpjos1QZl8fvXaF
GcDOqC9lrIxnmSydkMWoTerI2a/7yZiyQFpUyDHC2BPMNmRMEKWLywllVrDaTOzq
HAjfozO4S3zSifRySz3nxcfMXqwv8twtf8qSkYhoHBdcuQ/T3mTdoGzNsqIrH3Uf
8kG02bLEthDLIsMWHb2mod02+BYzm0BKvw0PiTxKF3udAVK/x83DIjJafqQXiNgr
gnuBtjAQX888kJPanp4f6a8brbDWm/+vq3uiFkMFRy4WP7Ycxfj7/7i14K+Hj/aN
IrLX8nmWMqaP7epIVGfw2mLjD2tAkeRmlxqMNxOu0El0xA5DO2G4BXO4ownOhWVF
bzi+j12aTJRqp6o246SvfoqaXGcW0am1nE+RL1pqtLuLUGRInOS28G7Ne9UAtpg0
7MjJZXyeQAmb21G2UAVqiF3JJdr87CjGOY6rAAKe/O8KWTYE1t/nca7NdSYFqOX2
N2+cqdnIGeA4oSmWqjS2xIVyxOgChHmG5XV9SFeeLXfzjHFl00yiw+580VIbLtHO
U0tuJRRiNQmZvPLlh1vqGLvzIGuyCd6/PonnbFZRoCtxRnG1/YVbXI8TSoSxHRnc
mCcjO8DRaSBvCWl7sA2h//57+4Ri8csx+Ml+doUxKiFrS9lVekvwYjKVNmFULJZw
IpGnGbw4HX50CiPgQPvXCXzGFPNTvrz1+ryT5p4l6BRoDQeplumlwftdCf8MVEaN
d9aUKo9xnaYegDb6rJT1PZfvtuj7hSOo/VnO0sl0zIDo9+B91ZRPemSxDEg2SJ3W
FL5UGK+VxTY7pAuvTOEwYpz2q+ITTGuyq6zDC1vYDuCid/Hf/UvXZITU20VxhUxn
/fGxyPZTKny00tENEUY6PHKF1giZklwjldlVjjSdC3cyvk6rxxEp8Qy5rQ/qy+o+
75BcVQwvMhdPs2bfcmK2HKnBYl4OX+8kW+2p04mONqiXk/6L9W7ldnTAonAUyxWb
k7ryxMaI2tq3MFwqbFhOf1v2wfcDWvlRHvwsTwQ+XvPbInoTFFuJ7Sbb+OTY5+8b
0lrabMObHVoQPKWNpE/xYzTjxgqj0aRpWYe9Qw6WT0dXT/21JfEeHftCm6RKA8YG
DoYBqlf6tqRj8Z6suLuePvrv8kJpDiY8PIwrzzetul4szD0X08WvAiA74+Txt2eN
Q3hdTwNH3lr0uqL/LunLBcHnoZIn2bTEL9vvffQYOP+9/fjLe3wqu2Vd6QxfdrIJ
RLtdtDcQ5PUbAyJZw59lw37Hsa5dC0R70rXh1uAzYAG3IIyVavGqgy5GOm8X0Tuj
gBR9SfyDgjUBQm6NJzf8+s2A4yzY0vNFbBL2NB/4t/c9iGeTXEn/3SvjTno6N2Z2
WlCm3a1jnP6cZuGWs0i/W1dpHe8De4FQ+WWxWm31G87q1Ez6E17IiKwfjVuOwnSt
xLByoaxiy+6BhJqp+V0/ibmon55QKUJqkWkfXsQGzMVUDVetNwai/OnTnS2Un3vM
IT7/L4Z5iheRW4ZixYIVipG7YDdAxV/gX+pB2sCLfLTwvQEfsVEEuPuTtzC8bbRE
y+Z5dUIBzY7R+T87Xzw3xsNeLulzFkDPfMHfZTViFejUIjwXsnQJ4k9mMjwGtouf
u7blTJLYYpU8+G9O03cCbaVrfaUaXdnBAbmkW23O8SaHRlOlybAe2eC+gkr3qgZR
91WzfDPyz2DFbBGGH76NPvGQUWeQkkIzEuWPUfzDXfliH9HYMpxb20twnQ46djnB
tDn/uvYSlQwuXfK6ydP5ET835sDU0MeA6zjqrPkbe4gHbTPj7MxKpiY+/Lq688XZ
XjSPfK73etjPrjp4ZHaP1ydcM+YnMqa2/uc2G5n+gvc8rI/OnQmDprIyLb/FJOpr
ICBTPMYoNs+dUK1l+MrCPq7i0YL4W4KmoasztKt3X7WGxU50vmEFxM/6AiRtJYLW
T8Rk4HOUtoMocSIRkbyT8iE2DYbu3gcUoWWW3dlyzPK3DYsEypfII7NPHmypfKOx
DyU7zM7E7LFwejHxdWrXg8sDuvdLJoI5uqhwQEIXnbYKPdwBDOPLHqctTM3PMNGV
i+VH+279IKcU0h124RKEHV/zJQpg7Tc5BaYEyjeTCt9kIdJzVB/OZHRGT5+Jq0BD
PDXgQ8GlZK/2a1kVXuDJLI503903Ew9TGZS6FyMg9b8ggwhNirVqFRYvr7DoL0kf
Yy96wYRrxwyf/tbefatENsMeJbANvcyfiy8BWRwafz96jdxDH/KMDTCfJzhKQ6g5
7Lo/BGKwUbUGoCCKykCq7MZaNmvYXfOMpkgv3WCnMik+IxljNcmRwXI1/4wuiMie
tKiGd9vvU0X/MSt/KDgJ5hvocsCi54BDEw30VB58Z0L+GwegtHENsuCIWvfmtwlA
2YvO3UOBAJHzYvevPf8dQf3RR0c6IDH9OzLuZ91c6pZ99PgLryTTGLaWBTFC42Y8
FXsW1Oqynu9JBIoT/Lg2nmokQsiX1lsMoRIzZp6jRy+8/3k+8lHBos/x8hmJVZxL
gbWbnGwJoaRzOO4+8SGHrh0VPL6knfq3KGjg5TxcdkBKJZHelQ937xlvSdK31DH1
7eMkdvE8aCvtQC8m5VBV8WR9rtyP4mCPtOHqPNiEoxwuTpXMyB5Ktf5uvjOFV9zB
BQ2/qoNlAa2C2e0i6rCaEYs1JZirMIBlu+v0gp9TIcAvbQqXLSfEr8Yq/an4WjOF
UJqiMw/Ky0FQM9vAuKDWfcZXaZNwvViCkooyEA/s9MoB4gMwrxP3rCs9QJVOaQvo
VJ4C+v97YWTf6jmy4CabxS+UZTTc5cPY4fWTP0+DDIGphw4VRq5JuWG3jQz1ogsY
Y8hW8dhgl8UmomM7ta7AuLZIUZoxoFJCFK5M22jdDU3KyHHyxF8YLxH6LvrX/vOW
gKWCP2nUdfWSbPued2Znr20XmmjUS65PIL9Lbox6O2gRsTqLFAbK9LButFICYt5m
JdzfH3MrCfpbhq93hjLRwNn2jXf8fzvMtReaUqSpprLExJNb7RU5a0QGOYhwSMuc
hFd1weoQT/b/dG1WdL8iv4n/zSvtg3aCIWOSf9rnYd2yBjZIGCNJqiJni3geKaOk
543lzNlyDM9/Wzw7wWB2uUJLCuD2FUlD9+yunrQwzb7fIzsey2PXrTSWeKMsM9+1
ZWljXSap4KnVNXydbWWOzTtpflpzV1R//Qh02RgX+5UTK++XGcUaf/+/twJRy+pT
AWgWYthQyW4OgqwsKzrofbDK3G4rzHeTBaV/ehveH0Ka52RosmpQFRgCrgnXXzpf
a3vnT1dP9pxd0tkMYPyPUirUP4WKa6RtChN8b+GA3Uf2k8EYzgZT1fcWZ9fGU2pN
8egQugV0VXtvAcilZunW/JCEB5thnFCZa5AGZvaBsmn4YP2ZMkjUqmVny4BRbuos
5DjWq1EULUrL2A5HIzkRJPudQuwYIVCo1lFdTUA1QZ21h6I8RgUfSTiE7QBOFcC0
IHatqF0H//VyjXF+DiPZz2eQ+9qF8PRDr62MZhN8VMQA16ppl1bHIu84tfueNIe1
2IJeJhBqv/23GEuPqHTIQdCGDLQ2TDR8NjQkV83sXND0ExHSExtw6YzBEECViY6P
ReW19UYUcQF9M4EsBzSJo34RnkXqAHXJ4etlHX7lmwDetAHJ1seg6SW6dk8eR8WN
t5GPNUo6u3vvs+WtS4bMT9X9YKtbp4iOWVeY6pG5fwI/QvXXt7bnI7qkwMYOsO+W
13fyKcFq0OpYth1F5/MQw0OeHaO+VWzHKLbmNXlz8HK/ozbVV1gzdzUGC4ySkLcN
1x7zo+qpTkLxT4zhZ739zwWHi5hbupbs7eYJjMsbiMca3oR/dMrlyb0W0J6q/+EN
QAoAL9Qm0MU3G3XAi7dEXxfFTUn5AT1MM3bwq93t0C8/d8iVTxALUb35EKRW1SoL
GbLJJx4dr2rQAtfagJUJzgdbQHRq1E1MvD5vlXPlhDly5xCzupyji3RRaKG1L2zb
pvYlLT38N5yf/pdDZZiTOr3UCR8ofwfaXmtwvqmr8XCh0ORWOjKpZnPm/nr3aQU6
EFdWsC6y8jV09uviLECda6cwPJ4aEeaL8jW9TxRu5gjp6itRxw9NLbuOvfr1xPTg
Uby4GQjue8smHsohAZqM8C2zHfS4n3ioE+jRznH9k4Fxz5XT5JCnQKKgzFPMU7pR
H/z8OUTt6Jgg1O76EKqv5vf15AJaifY+rwSUFbb+UcU5Vxbr+6IltYwY0k9IxzsR
hfF9WO192VgEKf1JKaB85c/T+0ydua8vUB3VvNFhXBYw5z5P+A71UBY51IZ7rYir
fWBA5ZhlQlqD5FadXxjV09rQDziSYQl9bYkvZliVFRNCCnBTaSd35CiUGy3QL9ul
bis5gs1IyDAPPrc9rkhToltgVFeTF+FZMDBhw2X/JMRbAzt908wcoP1Djuis7mkz
9PX8L+7oAuzWDlc73OYzZ4vynNy9+nJTy98fM5GR2w36Jlitum9ekrEdZbyRIP9g
tE1mynie5E9s3F5zQlkG7tv5upJ3Wm3XpIgpLZYvym6tAyKG3iOct2pER0cY6neQ
dbvfOGSG5GaxjzZ4bFHO8gDIWeGsYCQxMudwGyKlkAIQyV4dJtzcI2wf3gcdHZ2X
J3PL0+kqpwVIC80wE8qK1+dnzI3QEEU+JNtJu+3/aCUIZvUo/Nyb2/6nWzHBxXwq
dQKIAfpE2F9vbQ+5UfSfeqijEGHy3zG1zjFAWzNCjLEFtcDVqFghsYYEvjoStm/1
iWis61DjWsFiG9wEBC6Kjl9Eyxvgf26JjUgwlDmYFe01FUH5XRMUvD1h5aVlgGaj
5YpFytl7zmFPhK5LirRs9IS6weptljrEoWPHiVKDevOTPoipm2dXgw84oFrCxxst
aVG2C+OYsu4wkognbdogWjmnAiHAsZFut5ar6cscGOcoiufsghhMx9Sn2XlPxML6
rWkrqLfGHUnCSercHX2SBckcwojNBW+GgwUyCAXxXHHSmw3GmN2VpIzttbFwKnrS
UX1ZL0+LS1PSgm9S25pv7l9SI7nIsx+PiUEu6bHvDU7p3Ma/kVSKPvnOwP5Ptj8H
TU87fHfcOeRjLqYoyZ8qFNHquEhPeB2IifYYiQrlE6jpDaND8xjf9okG8cWKVcpd
7lwXUUJ2OeGOehmuPv7OkfRGakJfZ8d3+Vs5tBtqmJKSqRX8AUVxxZSOFlFNT9Bf
AQBuwFne9ybY9xXtZn1BPeDAn3gGH2GQJLx+AE4G9crRCgjnkZvnwzXf39MlsYSC
ckeqgufgJRCw1KSfCdrRqY6mhHO5Nyi4Xw1KX+YlCuxsgrvKeeFnOuaIBUIcWo1S
D2kvHffFYU7CY/X5Q6IKZ3JJUxfjeay8111Wb+o2pUynQlbNrZ5T677Ot9LdbY9V
2UBC280aBc4XOMq2lbKmryGsafwam2ZF5LAiP9RPaq/TxEjP6i7uwO4ltmCXQUab
kcpVXkmifxOrc5ihbqHQ+dgqyaKB2UKu2h52ezVQsAot9DXTYxUsxOTAc5CKH0+/
7bEMy5PqXiYa6doYcBIcHj49H5sqCjc2nICT+C7KWBQnOqxcRSuJVAi9CZv9AUnx
3P7M7yiReNCRdE8G48FK45bTzWk4WyE0VdmGiaz98Hl7H/HgWixNZyWZDRjBz4gj
0YitlR/aut9KF/8Au88jDdPM5fJnjK/WIi1YmAbg25v5bvSM15CrF5VxcHJBSqMR
emtVWX+SEWLUHDqVaP+Iy2+6rRrHEeY+H8JitFWpJfQA2rcobjHBVKOIEw2eHJqv
Xg/19bZ2HJXOfORTq8kPkF86g+TmUkKEyilQ9zpMUXNXlJIaPRuUk3dzrZabOBL5
dO3b+koFA9zgEywbHaNDKbe1GxAK+p4gzcHIhlXgxP6uQZMEN+GaXpMM0HnSlleG
hg8Iyq9ZmoB8KYMPfhWmEC9kwlKUzdfzCD4g7YiQ9VQ741q6Vuogw9+3KKqp/qvl
kg4Y5dCzj9bhdDtfIxxIj4s+LSaWr1Pf9uPMavp255usUSKWrw3SrE7mm95o3o6d
W1Pno50rMg8PGVIPy+2gYhLyNfMFqXtXwz99lopeNYlDhQed5Oiu/nGNPSjJ44ug
Z4dg133XD+nK2RF85X3AwNBeegpkLWP2Ke3BTla8zWIZMNOBmgUEOuUqt+8YsgJ6
O6sbPhNalcTkK9VP/PlwqkA/TrVTYEjmVfZ5M6eCxPEUub6wxNS+X1Rgf+5iYQDn
FdrTapF6SBIUu8KX+fzl6EjGthpR8JV012dLVe7sTEnugRiBs9GW9RmQfEB0sNsd
NqkZcIifVk2heYTkWotukJtAGyYY9h6hx7noAxs6h8+8q1xtJotTO3uhcLqsTck/
W0pyqEdoV+SqrnErIjZWZ3bSQqnKLlYAOu6zdg5M8Pfi+FhTFfo65AfPpCyPyY1d
nqRolvePMEe52WMCHihOOrcJN3RW8Q7F9tzn1WXH81euAYXhliyG1JWGjyu3N0sr
SiEfersjmS9j+YXdbXevLd0ftfUnxL8M12PaO0wL0pVqVCBI9+cmdtEOZYXQIBJp
mEPjevA0lbGPVO+QfvS2YdQY6O76HRvTQx2kej0V+kzmg6+5l2gxW6Bxnx5xkINZ
R+z5RXfZbUj4SH5C54tQWhyYYNtKa7EkuHY4JYCQwaV0oJMec5IqBs8Jz/2Qua5B
uOuP7naJ99Gc529eEci/kezg0C1kwruXixOdcz4TGkSL7aa5XA5gqPtacapHBCas
UxxxaXqWV4xXLm7FBbY6IIG0I7KXZUEWQ3+VtCyAW/oHzYKxrugyHxEqmIRAtRw7
37sYhxe5exfsgr5tj3dPzSrCL0fheFhlGiNgCyq2gYUUtCugzTfTEuwXTVP0ufuh
Ld1lLWaeLGWaTJcxkyBGdeMsu6eXC4G3+8AkSJpPbY46kYBOBKPsCKMSBrRFe+Tv
Pbbjlkmsh45r9ZwtGLkxskjZcI4OrrWK87usKXoTaABXg7Fac2+kjxOn3qhN2RVn
i6xTWHZwBClnkqDjyzI3A8mbjN4I622Se4EhzNu2iwggR5273ekB/FiZsknloV3l
K5uVQpegxhZggJwLwD07M46uja5C/9gvhz/Qo7kHTyrOlcoptUvhD/AmokMpx/4H
381lIxXCw2LZzfX+FxvbOW3GAwLcOAfQu+waRyLQRQtRyo15VzQWBwcKbvR5MGHJ
umY+Ji7MG2BcxZGrq/1yA5wmBC2imzCSl4BitbJVagmEdfE77ownzCLi++ctvpbn
S+JNMufO6pgvV//J13gJsXlS7hNjChCrozQrjMwyKgr7nLLvzhh3a2BpAPLTLGEy
7umkZ4ttczwiKq3ANMQr46/XnNEGaHVkWSr5gy+50aIooMHsclz2UDUKmxmBz+OO
4fHbKyGPYrbmlx+ALqTcV3Wjd0EuFyBRtK5ylQtNrGmtMafRUh4gTtl6g9SQJja2
t6hX/jhxGh3oMSbeLtqteAdbLTbBpK4VTEycBfk2yxW/a1ujdVs3DyyjL4ceTS2A
ogu0iAbzkA8mWsSMKaUfRzj/cLr7P5QJ278ST6QrEdLvfLdtcYkm4r6MwnKuWBNu
J+Y2PmxJPGZo6tuj8yztEceLBDPOYa2curLjKAoT4a1I3u/QiWV7RQnYI6+zSXVv
NxfumiAD+QHLksb9vVsPdg5w/DiZwwlEpqKADPjEIe21r0bfeorHkFTSCgLctT6S
mSliR0qMC90ZJAFtWuZWOdnT7l0/Jlw0z6W/QTjqqdx4y/h6OZzFu1vxtmrfOsXY
iYiMFE6FNygvWMSDW3lGmxenGg/wdVMRfa5q68lVhY8Ywre/BDKV4IGECuQ79oyz
MFPLUu+Jjvf0xVmzIKCMzK9yGk3xW/ip0+aHErmuyNgCWdiVguOl7J5rslzkWBj8
VGlqJbjGGKqiQEg6YEa14lYIAFYlCufwjzrtOSokb9Y=
`protect END_PROTECTED
