module tile_router_v1_00_a_output_arbiter(clk,rst,enable,requests,requests_accept,select_valid,select,select_oh);
input clk;
input rst;
input enable;
input [7:0] requests;
output reg  select_valid;
output reg [2:0] select;
output reg [7:0] select_oh;
output     [7:0] requests_accept;

reg [2:0] select_c;
reg [7:0] select_oh_c;
reg [7:0] tie;
reg [7:0] tie_c;

always@(posedge clk)
begin
	if (rst)
	begin
		select_valid <= 1'b0;
	end
	else
	begin
		if (enable)
		begin
			select_valid <= |requests;
		end
		else
		begin
			select_valid <= 1'b0;
		end
	end
end

always @(posedge clk)
begin
	if (rst)
	begin
		tie <= 8'b00000001;
		select_oh <= 8'b0;
		select <= 3'b0;
	end
	else
	begin
		if (enable)
		begin
			tie 		<= tie_c;
			select_oh 	<= select_oh_c;
			select 		<= select_c;
		end
	end
end

assign requests_accept = select_oh_c;

always@*
begin
	
	(* full_case *)case({tie,requests})
		16'b10000000_00000000 : begin select_oh_c <= 8'b00000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_00000000 : begin select_oh_c <= 8'b00000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00100000_00000000 : begin select_oh_c <= 8'b00000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00010000_00000000 : begin select_oh_c <= 8'b00000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00001000_00000000 : begin select_oh_c <= 8'b00000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000100_00000000 : begin select_oh_c <= 8'b00000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_00000000 : begin select_oh_c <= 8'b00000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_00000000 : begin select_oh_c <= 8'b00000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_00000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b01000000_00000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00100000_00000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00010000_00000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00001000_00000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_00000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_00000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b01000000_00000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00100000_00000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00010000_00000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_00000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_00000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b10000000_00000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b01000000_00000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00100000_00000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00010000_00000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_00000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_00000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00000011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b01000000_00000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00100000_00000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_00000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_00000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000001_00000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b10000000_00000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b01000000_00000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00100000_00000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_00000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_00000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00000101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00000101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b01000000_00000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00100000_00000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_00000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_00000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00000110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b10000000_00000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b01000000_00000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00100000_00000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_00000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_00000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00000111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00000111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b01000000_00001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_00001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_00001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000010_00001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000001_00001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b10000000_00001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b01000000_00001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_00001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_00001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_00001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b01000000_00001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_00001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_00001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00001010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00001010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b10000000_00001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b01000000_00001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_00001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_00001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00001011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00001011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00001011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b01000000_00001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_00001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_00001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00001100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000001_00001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b10000000_00001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b01000000_00001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_00001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_00001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00001101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00001101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00001101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b01000000_00001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_00001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_00001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00001110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00001110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b10000000_00001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b01000000_00001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_00001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_00001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00001111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00001111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00001111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00000100_00010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00000010_00010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00000001_00010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b10000000_00010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_00010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_00010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_00010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b10000000_00010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_00010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00010011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00010100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00010100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00000001_00010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b10000000_00010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00010101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00010101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00010101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00010101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00010110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00010110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00010110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b10000000_00010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00010111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00010111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00010111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00010111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00011000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00000010_00011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00000001_00011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b10000000_00011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00011001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_00011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00011010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00011010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00011010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b10000000_00011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00011011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00011011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00011011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00011011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00011100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00011100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00000001_00011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b10000000_00011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00011101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00011101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00011101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00011101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00011110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00011110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00011110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b10000000_00011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b01000000_00011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_00011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_00011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00011111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00011111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00011111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00011111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00001000_00100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000100_00100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000010_00100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000001_00100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00100001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00100001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00100001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00001000_00100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_00100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_00100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00100010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00100010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00100010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_00100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_00100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00100010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00100011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00100011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00100011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_00100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_00100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00100011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00100100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00100100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00100100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_00100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00100100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000001_00100100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00100101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00100101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00100101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_00100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00100101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00100101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00100110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00100110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00100110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_00100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00100110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00100110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00100111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00100111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00100111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_00100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00100111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00100111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00101000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00101000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000010_00101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000001_00101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00101001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00101001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00101001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00101001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00101001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_00101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00101010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00101010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00101010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00101010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00101010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00101010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00101010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00101010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00101011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00101011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00101011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00101011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00101011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00101011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00101011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00101011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00101100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00101100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00101100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00101100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00101100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00101100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00101100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000001_00101100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00101101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00101101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00101101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00101101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00101101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00101101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00101101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00101101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00101110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00101110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00101110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00101110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00101110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00101110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00101110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00101110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00101111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00101111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00101111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00101111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_00101111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00101111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00101111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00101111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00110000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000100_00110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000010_00110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000001_00110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00110001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00110001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00110001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00110001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_00110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_00110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00110010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00110010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00110010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00110010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_00110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00110010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00110011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00110011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00110011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00110011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_00110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00110011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00110100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00110100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00110100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00110100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00110100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00110100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00110100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000001_00110100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00110101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00110101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00110101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00110101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00110101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00110101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00110101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00110101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00110110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00110110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00110110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00110110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00110110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00110110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00110110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00110110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00110111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00110111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00110111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00110111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00110111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_00110111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00110111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00110111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00111000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00111000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000010_00111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000001_00111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00111001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00111001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00111001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00111001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00111001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_00111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00111010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00111010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00111010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00111010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00111010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00111010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00111010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00111010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00111011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00111011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00111011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00111011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00111011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00111011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_00111011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00111011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00111100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00111100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00111100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00111100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00111100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00111100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00111100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00000001_00111100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00111101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00111101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00111101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00111101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00111101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00111101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00111101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_00111101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_00111110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00111110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00111110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00111110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00111110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00111110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00111110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00111110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b10000000_00111111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b01000000_00111111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_00111111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_00111111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_00111111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_00111111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_00111111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_00111111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01000000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01000000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01000000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00010000_01000000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00001000_01000000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000100_01000000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000010_01000000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01000000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01000001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01000001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00010000_01000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00001000_01000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_01000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_01000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01000010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01000010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00010000_01000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_01000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_01000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01000010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01000011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01000011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00010000_01000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_01000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_01000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01000011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01000100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01000100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_01000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_01000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01000100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01000100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01000101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01000101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_01000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_01000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01000101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01000101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01000110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01000110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_01000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_01000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01000110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01000110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01000111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01000111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_01000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_01000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01000111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01000111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01001000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01001000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_01001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01001000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000010_01001000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01001000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01001001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01001001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_01001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_01001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01001010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01001010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_01001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01001010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01001010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01001010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01001011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01001011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_01001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01001011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01001011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01001011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01001100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01001100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_01001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01001100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01001100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01001100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01001101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01001101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_01001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01001101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01001101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01001101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01001110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01001110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_01001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01001110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01001110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01001110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01001111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01001111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_01001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01001111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01001111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01001111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01010000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01010000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01010000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000100_01010000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000010_01010000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01010000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01010001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01010001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_01010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_01010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01010010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01010010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_01010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01010010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01010011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01010011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_01010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01010011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01010100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01010100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01010100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01010100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01010100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01010100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01010101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01010101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01010101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01010101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01010101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01010101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01010110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01010110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01010110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01010110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01010110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01010110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01010111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01010111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01010111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01010111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01010111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01010111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01011000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01011000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01011000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01011000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000010_01011000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01011000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01011001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01011001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01011001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_01011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01011010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01011010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01011010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01011010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01011010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01011010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01011011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01011011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01011011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01011011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01011011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01011011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01011100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01011100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01011100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01011100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01011100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01011100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01011101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01011101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01011101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01011101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01011101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01011101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01011110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01011110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01011110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01011110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01011110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01011110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01011111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01011111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_01011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01011111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01011111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01011111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01011111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01100000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01100000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01100000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00001000_01100000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000100_01100000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000010_01100000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01100000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01100001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01100001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01100001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00001000_01100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_01100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_01100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01100010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01100010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01100010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_01100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_01100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01100010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01100011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01100011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01100011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_01100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_01100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01100011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01100100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01100100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01100100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_01100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01100100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01100100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01100101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01100101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01100101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_01100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01100101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01100101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01100110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01100110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01100110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_01100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01100110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01100110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01100111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01100111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01100111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_01100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01100111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01100111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01101000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01101000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01101000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01101000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01101000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000010_01101000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01101000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01101001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01101001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01101001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01101001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01101001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_01101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01101010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01101010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01101010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01101010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01101010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01101010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01101010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01101010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01101011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01101011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01101011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01101011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01101011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01101011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01101011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01101011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01101100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01101100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01101100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01101100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01101100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01101100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01101100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01101100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01101101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01101101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01101101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01101101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01101101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01101101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01101101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01101101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01101110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01101110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01101110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01101110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01101110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01101110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01101110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01101110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01101111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01101111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01101111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01101111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_01101111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01101111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01101111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01101111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01110000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01110000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01110000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01110000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000100_01110000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000010_01110000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01110000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01110001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01110001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01110001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01110001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_01110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_01110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01110010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01110010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01110010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01110010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_01110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01110010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01110011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01110011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01110011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01110011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_01110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01110011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01110100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01110100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01110100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01110100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01110100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01110100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01110100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01110100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01110101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01110101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01110101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01110101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01110101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01110101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01110101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01110101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01110110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01110110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01110110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01110110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01110110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01110110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01110110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01110110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01110111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01110111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01110111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01110111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01110111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_01110111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01110111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01110111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01111000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01111000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01111000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01111000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01111000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000010_01111000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01111000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01111001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01111001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01111001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01111001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01111001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_01111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01111010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01111010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01111010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01111010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01111010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01111010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01111010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01111010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01111011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01111011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01111011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01111011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01111011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01111011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_01111011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01111011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01111100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01111100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01111100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01111100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01111100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01111100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01111100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00000001_01111100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01111101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01111101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01111101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01111101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01111101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01111101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01111101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_01111101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_01111110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01111110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01111110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01111110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01111110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01111110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01111110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01111110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b10000000_01111111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b01000000_01111111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_01111111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_01111111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_01111111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_01111111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_01111111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_01111111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00100000_10000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00010000_10000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00001000_10000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000100_10000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_10000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10000001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00100000_10000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00010000_10000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00001000_10000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_10000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_10000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10000010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00100000_10000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00010000_10000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_10000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_10000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10000010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10000011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00100000_10000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00010000_10000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_10000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_10000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10000011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10000100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00100000_10000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_10000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_10000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10000100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10000100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10000101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00100000_10000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_10000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_10000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10000101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10000101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10000110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00100000_10000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_10000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_10000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10000110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10000110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10000111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00100000_10000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_10000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_10000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10000111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10000111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10001000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_10001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_10001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10001000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_10001000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10001000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10001001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_10001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_10001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_10001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10001010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_10001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_10001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10001010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10001010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10001010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10001011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_10001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_10001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10001011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10001011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10001011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10001100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_10001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_10001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10001100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10001100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10001100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10001101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_10001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_10001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10001101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10001101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10001101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10001110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_10001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_10001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10001110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10001110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10001110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10001111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00100000_10001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_10001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10001111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10001111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10001111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000100_10010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_10010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10010001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_10010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_10010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10010010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_10010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10010010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10010011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_10010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10010011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10010100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10010100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10010100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10010100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10010100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10010101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10010101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10010101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10010101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10010101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10010110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10010110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10010110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10010110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10010110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10010111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10010111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10010111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10010111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10010111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10011000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10011000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10011000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_10011000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10011000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10011001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10011001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_10011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10011010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10011010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10011010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10011010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10011010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10011011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10011011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10011011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10011011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10011011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10011100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10011100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10011100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10011100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10011100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10011101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10011101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10011101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10011101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10011101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10011110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10011110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10011110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10011110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10011110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10011111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00100000_10011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_10011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10011111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10011111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10011111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10011111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00001000_10100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000100_10100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_10100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10100001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10100001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10100001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00001000_10100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_10100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_10100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10100010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10100010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10100010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_10100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_10100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10100010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10100011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10100011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10100011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_10100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_10100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10100011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10100100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10100100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10100100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_10100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10100100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10100100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10100101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10100101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10100101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_10100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10100101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10100101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10100110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10100110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10100110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_10100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10100110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10100110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10100111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10100111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10100111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_10100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10100111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10100111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10101000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10101000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10101000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10101000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_10101000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10101000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10101001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10101001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10101001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10101001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10101001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_10101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10101010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10101010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10101010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10101010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10101010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10101010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10101010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10101010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10101011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10101011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10101011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10101011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10101011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10101011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10101011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10101011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10101100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10101100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10101100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10101100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10101100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10101100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10101100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10101100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10101101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10101101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10101101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10101101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10101101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10101101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10101101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10101101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10101110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10101110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10101110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10101110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10101110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10101110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10101110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10101110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10101111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10101111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10101111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10101111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_10101111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10101111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10101111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10101111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10110000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000100_10110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_10110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10110001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10110001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10110001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10110001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_10110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_10110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10110010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10110010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10110010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10110010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_10110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10110010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10110011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10110011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10110011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10110011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_10110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10110011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10110100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10110100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10110100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10110100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10110100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10110100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10110100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10110100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10110101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10110101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10110101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10110101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10110101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10110101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10110101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10110101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10110110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10110110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10110110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10110110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10110110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10110110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10110110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10110110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10110111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10110111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10110111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10110111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10110111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_10110111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10110111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10110111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10111000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10111000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10111000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10111000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_10111000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10111000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10111001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10111001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10111001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10111001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10111001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_10111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10111010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10111010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10111010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10111010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10111010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10111010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10111010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10111010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10111011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10111011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10111011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10111011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10111011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10111011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_10111011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10111011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10111100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10111100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10111100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10111100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10111100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10111100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10111100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_10111100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10111101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10111101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10111101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10111101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10111101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10111101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10111101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_10111101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_10111110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10111110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10111110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10111110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10111110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10111110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10111110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10111110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_10111111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_10111111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00100000_10111111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_10111111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_10111111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_10111111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_10111111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_10111111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11000000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00010000_11000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00001000_11000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000100_11000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_11000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11000000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11000001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11000001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00010000_11000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00001000_11000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_11000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_11000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11000001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11000010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11000010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00010000_11000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_11000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_11000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11000010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11000010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11000011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11000011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00010000_11000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_11000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_11000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11000011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11000011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11000100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11000100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_11000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_11000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11000100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11000100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11000100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11000101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11000101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_11000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_11000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11000101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11000101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11000101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11000110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11000110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_11000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_11000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11000110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11000110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11000110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11000111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11000111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00010000_11000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_11000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11000111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11000111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11000111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11001000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11001000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_11001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11001000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11001000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_11001000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11001000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11001001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11001001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_11001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11001001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_11001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11001001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11001010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11001010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_11001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11001010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11001010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11001010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11001010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11001011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11001011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_11001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11001011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11001011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11001011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11001011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11001100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11001100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_11001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11001100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11001100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11001100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11001100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11001101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11001101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_11001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11001101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11001101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11001101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11001101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11001110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11001110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_11001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11001110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11001110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11001110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11001110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11001111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11001111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00010000_11001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11001111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11001111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11001111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11001111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11010000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11010000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000100_11010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_11010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11010000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11010001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11010001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11010001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_11010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_11010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11010001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11010010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11010010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11010010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_11010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11010010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11010010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11010011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11010011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11010011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_11010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11010011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11010011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11010100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11010100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11010100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11010100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11010100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11010100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11010100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11010101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11010101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11010101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11010101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11010101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11010101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11010101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11010110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11010110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11010110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11010110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11010110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11010110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11010110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11010111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11010111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11010111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11010111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11010111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11010111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11010111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11011000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11011000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11011000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11011000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11011000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_11011000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11011000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11011001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11011001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11011001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11011001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_11011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11011001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11011010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11011010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11011010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11011010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11011010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11011010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11011010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11011011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11011011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11011011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11011011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11011011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11011011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11011011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11011100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11011100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11011100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11011100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11011100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11011100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11011100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11011101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11011101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11011101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11011101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11011101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11011101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11011101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11011110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11011110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11011110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11011110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11011110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11011110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11011110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11011111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11011111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00010000_11011111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11011111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11011111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11011111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11011111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11100000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11100000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00001000_11100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000100_11100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_11100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11100000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11100001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11100001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11100001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00001000_11100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_11100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_11100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11100001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11100010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11100010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11100010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_11100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_11100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11100010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11100010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11100011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11100011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11100011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00001000_11100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_11100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11100011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11100011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11100100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11100100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11100100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_11100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11100100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11100100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11100100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11100101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11100101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11100101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_11100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11100101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11100101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11100101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11100110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11100110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11100110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_11100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11100110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11100110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11100110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11100111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11100111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11100111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00001000_11100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11100111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11100111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11100111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11101000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11101000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11101000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11101000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11101000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11101000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_11101000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11101000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11101001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11101001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11101001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11101001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11101001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_11101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11101001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11101010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11101010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11101010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11101010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11101010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11101010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11101010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11101010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11101011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11101011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11101011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11101011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11101011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11101011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11101011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11101011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11101100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11101100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11101100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11101100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11101100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11101100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11101100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11101100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11101101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11101101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11101101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11101101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11101101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11101101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11101101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11101101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11101110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11101110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11101110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11101110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11101110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11101110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11101110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11101110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11101111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11101111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11101111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11101111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00001000_11101111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11101111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11101111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11101111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11110000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11110000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11110000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000100_11110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_11110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11110000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11110001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11110001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11110001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11110001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000100_11110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_11110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11110001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11110010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11110010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11110010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11110010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_11110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11110010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11110010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11110011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11110011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11110011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11110011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000100_11110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11110011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11110011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11110100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11110100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11110100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11110100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11110100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11110100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11110100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11110100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11110101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11110101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11110101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11110101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11110101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11110101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11110101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11110101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11110110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11110110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11110110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11110110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11110110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11110110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11110110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11110110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11110111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11110111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11110111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11110111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11110111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000100_11110111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11110111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11110111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11111000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11111000 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11111000 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11111000 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11111000 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11111000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000010_11111000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11111000 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11111001 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11111001 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11111001 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11111001 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11111001 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000010_11111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11111001 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11111010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11111010 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11111010 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11111010 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11111010 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11111010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11111010 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11111010 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11111011 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11111011 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11111011 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11111011 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11111011 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11111011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000010_11111011 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11111011 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11111100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11111100 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11111100 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11111100 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11111100 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11111100 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11111100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b00000001_11111100 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11111101 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11111101 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11111101 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11111101 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11111101 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11111101 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11111101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b00000001_11111101 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
		16'b10000000_11111110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11111110 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11111110 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11111110 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11111110 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11111110 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11111110 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11111110 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b10000000_11111111 : begin select_oh_c <= 8'b10000000; select_c <= 3'b111; tie_c <= 8'b01000000; end
		16'b01000000_11111111 : begin select_oh_c <= 8'b01000000; select_c <= 3'b110; tie_c <= 8'b00100000; end
		16'b00100000_11111111 : begin select_oh_c <= 8'b00100000; select_c <= 3'b101; tie_c <= 8'b00010000; end
		16'b00010000_11111111 : begin select_oh_c <= 8'b00010000; select_c <= 3'b100; tie_c <= 8'b00001000; end
		16'b00001000_11111111 : begin select_oh_c <= 8'b00001000; select_c <= 3'b011; tie_c <= 8'b00000100; end
		16'b00000100_11111111 : begin select_oh_c <= 8'b00000100; select_c <= 3'b010; tie_c <= 8'b00000010; end
		16'b00000010_11111111 : begin select_oh_c <= 8'b00000010; select_c <= 3'b001; tie_c <= 8'b00000001; end
		16'b00000001_11111111 : begin select_oh_c <= 8'b00000001; select_c <= 3'b000; tie_c <= 8'b10000000; end
	endcase
end
endmodule
