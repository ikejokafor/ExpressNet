`timescale 1ns / 1ns
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company:    
//        
// Engineer:  
//
// Create Date:    
// Design Name:    
// Module Name:    
// Project Name:  
// Target Devices:  
// Tool versions:
// Description:   
//                
//                
//
// Dependencies:  
//                
//                
//                
//    
// Revision:
//
// Additional Comments:
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
module clock_gen #(
    parameter C_PERIOD_BY_2 = 5
) (
    clk_out
);    
    // ----------------------------------------------------------------------------------------------------------------------------------------------
    // Inputs / Outputs
    // ----------------------------------------------------------------------------------------------------------------------------------------------
    output  clk_out;
    
    
    //-----------------------------------------------------------------------------------------------------------------------------------------------
    // Regs
    //-----------------------------------------------------------------------------------------------------------------------------------------------
    reg clk_out_r;
    
    
    // BEGIN Clock Gen logic ------------------------------------------------------------------------------------------------------------------------
    initial begin
		clk_out_r = 1;
	end   
    
    assign clk_out = clk_out_r;
  
    always@(*) begin
        #C_PERIOD_BY_2 clk_out_r <= ~clk_out_r;
    end
    // END Clock Gen logic --------------------------------------------------------------------------------------------------------------------------

    
endmodule



