library verilog;
use verilog.vl_types.all;
entity cnl_sc0_generator_sv_unit is
end cnl_sc0_generator_sv_unit;
