parameter  C_PACKET_WIDTH		= 66;
localparam C_DATAIN_WIDTH      = 18;
localparam C_WEIGHT_WIDTH_IN   = 32;
localparam C_WEIGHT_WIDTH      = C_WEIGHT_WIDTH_IN >> 1;
localparam C_A_INPUT_WIDTH     = 30;
localparam C_B_INPUT_WIDTH     = 18;

localparam C_P_OUTPUT_WIDTH   = 48;