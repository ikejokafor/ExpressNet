
`ifndef __TILE_ROUTER_V1_00_A_DEFINES__
`define __TILE_ROUTER_V1_00_A_DEFINES__

`define PACKET_WIDTH					66

`define SRC_DST_PE_WIDTH				2
`define SRC_DST_PE_LOW					0
`define SRC_DST_PE_HIGH					(`SRC_DST_PE_LOW + `SRC_DST_PE_WIDTH - 1)
`define SRC_DST_PE_FIELD				(`SRC_DST_PE_HIGH):(`SRC_DST_PE_LOW)

`define SRC_ADDRESS_WIDTH				6
`define SRC_ADDRESS_LOW					(`SRC_DST_PE_HIGH + 1)
`define SRC_ADDRESS_HIGH				(`SRC_ADDRESS_LOW + `SRC_ADDRESS_WIDTH - 1)
`define SRC_ADDRESS_FIELD				(`SRC_ADDRESS_HIGH):(`SRC_ADDRESS_LOW)
`define SRC_ADDRESS_X_WIDTH				3
`define SRC_ADDRESS_X_LOW				`SRC_ADDRESS_LOW
`define SRC_ADDRESS_X_HIGH				(`SRC_ADDRESS_X_LOW + `SRC_ADDRESS_X_WIDTH - 1)
`define SRC_ADDRESS_X_FIELD				(`SRC_ADDRESS_X_HIGH):(`SRC_ADDRESS_X_LOW)
`define SRC_ADDRESS_Y_WIDTH				3
`define SRC_ADDRESS_Y_LOW				(`SRC_ADDRESS_X_HIGH + 1)
`define SRC_ADDRESS_Y_HIGH				(`SRC_ADDRESS_Y_LOW + `SRC_ADDRESS_Y_WIDTH - 1)
`define SRC_ADDRESS_Y_FIELD				(`SRC_ADDRESS_Y_HIGH):(`SRC_ADDRESS_Y_LOW)

`define DST_ADDRESS_WIDTH				6
`define DST_ADDRESS_LOW					(`SRC_ADDRESS_HIGH + 1)
`define DST_ADDRESS_HIGH				(`DST_ADDRESS_LOW + `DST_ADDRESS_WIDTH - 1)
`define DST_ADDRESS_FIELD				(`DST_ADDRESS_HIGH):(`DST_ADDRESS_LOW)
`define DST_ADDRESS_X_WIDTH				3
`define DST_ADDRESS_X_LOW				`DST_ADDRESS_LOW
`define DST_ADDRESS_X_HIGH				(`DST_ADDRESS_X_LOW + `DST_ADDRESS_X_WIDTH - 1)
`define DST_ADDRESS_X_FIELD				(`DST_ADDRESS_X_HIGH):(`DST_ADDRESS_X_LOW)
`define DST_ADDRESS_Y_WIDTH				3
`define DST_ADDRESS_Y_LOW				(`DST_ADDRESS_X_HIGH + 1)
`define DST_ADDRESS_Y_HIGH				(`DST_ADDRESS_Y_LOW + `DST_ADDRESS_Y_WIDTH - 1)
`define DST_ADDRESS_Y_FIELD				(`DST_ADDRESS_Y_HIGH):(`DST_ADDRESS_Y_LOW)

`define TAG_WIDTH						4
`define	TAG_LOW							(`DST_ADDRESS_HIGH + 1)
`define TAG_HIGH						(`TAG_LOW + `TAG_WIDTH - 1)
`define TAG_FIELD						(`TAG_HIGH):(`TAG_LOW)

`define TYPE_WIDTH						2
`define TYPE_LOW						(`TAG_HIGH + 1)
`define TYPE_HIGH						(`TYPE_LOW + `TYPE_WIDTH - 1)
`define TYPE_FIELD						(`TYPE_HIGH):(`TYPE_LOW)

`define ADDRESS_WIDTH					14
`define	ADDRESS_LOW						(`TYPE_HIGH + 1)
`define ADDRESS_HIGH					(`ADDRESS_LOW + `ADDRESS_WIDTH - 1)
`define ADDRESS_FIELD					(`ADDRESS_HIGH):(`ADDRESS_LOW)

`define MESSAGE_CODE_WIDTH				6
`define MESSAGE_CODE_LOW				(`ADDRESS_HIGH + 1)
`define MESSAGE_CODE_HIGH				(`MESSAGE_CODE_LOW + `MESSAGE_CODE_WIDTH - 1)
`define MESSAGE_CODE_FIELD				(`MESSAGE_CODE_HIGH):(`MESSAGE_CODE_LOW)
`define MESSAGE_DATA_WIDTH				40
`define MESSAGE_DATA_LOW				(`MESSAGE_CODE_HIGH + 1)
`define MESSAGE_DATA_HIGH				(`MESSAGE_DATA_LOW + `MESSAGE_DATA_WIDTH - 1)
`define MESSAGE_DATA_FIELD				(`MESSAGE_DATA_HIGH):(`MESSAGE_DATA_LOW)

`define READ_REQ_HAAR_ADDRESS_ROW_WIDTH	7
`define READ_REQ_HAAR_ADDRESS_ROW_LOW	(`ADDRESS_LOW)
`define READ_REQ_HAAR_ADDRESS_ROW_HIGH	(`READ_REQ_HAAR_ADDRESS_ROW_LOW + `READ_REQ_HAAR_ADDRESS_ROW_WIDTH - 1)
`define READ_REQ_HAAR_ADDRESS_ROW_FIELD	(`READ_REQ_HAAR_ADDRESS_ROW_HIGH):(`READ_REQ_HAAR_ADDRESS_ROW_LOW)
`define READ_REQ_HAAR_ADDRESS_COL_WIDTH	7
`define READ_REQ_HAAR_ADDRESS_COL_LOW	(`READ_REQ_HAAR_ADDRESS_ROW_HIGH + 1)
`define READ_REQ_HAAR_ADDRESS_COL_HIGH	(`READ_REQ_HAAR_ADDRESS_COL_LOW + `READ_REQ_HAAR_ADDRESS_COL_WIDTH - 1)
`define READ_REQ_HAAR_ADDRESS_COL_FIELD	(`READ_REQ_HAAR_ADDRESS_COL_HIGH):(`READ_REQ_HAAR_ADDRESS_COL_LOW)
`define READ_REQ_HAAR_ENABLE_WIDTH		6
`define READ_REQ_HAAR_ENABLE_LOW		(`ADDRESS_HIGH + 1)
`define READ_REQ_HAAR_ENABLE_HIGH		(`READ_REQ_HAAR_ENABLE_LOW + `READ_REQ_HAAR_ENABLE_WIDTH - 1)
`define READ_REQ_HAAR_ENABLE_FIELD		(`READ_REQ_HAAR_ENABLE_HIGH):(`READ_REQ_HAAR_ENABLE_LOW)
`define READ_REQ_HAARX_FLAG				(`READ_REQ_HAAR_ENABLE_HIGH + 1)
`define READ_REQ_HAARY_FLAG				(`READ_REQ_HAARX_FLAG + 1)
`define READ_REQ_HAAR_INFO_WIDTH		(`READ_REQ_HAAR_ENABLE_WIDTH + 2)
`define READ_REQ_HAAR_INFO_LOW			(`READ_REQ_HAAR_ENABLE_LOW)
`define READ_REQ_HAAR_INFO_HIGH			(`READ_REQ_HAARY_FLAG)
`define READ_REQ_HAAR_INFO_FIELD		(`READ_REQ_HAAR_INFO_HIGH):(`READ_REQ_HAAR_INFO_LOW)
`define READ_REQ_HAAR_OFFSET_WIDTH		11
`define READ_REQ_HAAR_OFFSET_LOW		(`READ_REQ_HAAR_INFO_HIGH + 1)
`define READ_REQ_HAAR_OFFSET_HIGH		(`READ_REQ_HAAR_OFFSET_LOW + `READ_REQ_HAAR_OFFSET_WIDTH - 1)
`define READ_REQ_HAAR_OFFSET_FIELD		(`READ_REQ_HAAR_OFFSET_HIGH):(`READ_REQ_HAAR_OFFSET_LOW)
`define READ_REQ_RSVD_WIDTH				13
`define READ_REQ_RSVD_LOW				(`READ_REQ_HAAR_OFFSET_HIGH + 1)
`define READ_REQ_RSVD_HIGH				(`READ_REQ_RSVD_LOW + `READ_REQ_RSVD_WIDTH - 1)
`define READ_REQ_RSVD_FIELD				(`READ_REQ_RSVD_HIGH):(`READ_REQ_RSVD_LOW)

`define READ_REPLY_HAAR_ENABLE_WIDTH	6
`define READ_REPLY_HAAR_ENABLE_LOW		(`ADDRESS_HIGH + 1)
`define READ_REPLY_HAAR_ENABLE_HIGH		(`READ_REPLY_HAAR_ENABLE_LOW + `READ_REPLY_HAAR_ENABLE_WIDTH - 1)
`define READ_REPLY_HAAR_ENABLE_FIELD	(`READ_REPLY_HAAR_ENABLE_HIGH):(`READ_REPLY_HAAR_ENABLE_LOW)
`define READ_REPLY_HAARX_FLAG			(`READ_REPLY_HAAR_ENABLE_HIGH + 1)
`define READ_REPLY_HAARY_FLAG			(`READ_REPLY_HAARX_FLAG + 1)
`define READ_REPLY_HAAR_INFO_WIDTH		(`READ_REPLY_HAAR_ENABLE_WIDTH + 2)
`define READ_REPLY_HAAR_INFO_LOW		(`READ_REPLY_HAAR_ENABLE_LOW)
`define READ_REPLY_HAAR_INFO_HIGH		(`READ_REPLY_HAARY_FLAG)
`define READ_REPLY_HAAR_INFO_FIELD		(`READ_REPLY_HAAR_INFO_HIGH):(`READ_REPLY_HAAR_INFO_LOW)
`define READ_REPLY_RSVD_WIDTH			6
`define READ_REPLY_RSVD_LOW				(`READ_REPLY_HAAR_INFO_HIGH + 1)
`define READ_REPLY_RSVD_HIGH			(`READ_REPLY_RSVD_LOW + `READ_REPLY_RSVD_WIDTH - 1)
`define READ_REPLY_RSVD_FIELD			(`READ_REPLY_RSVD_HIGH):(`READ_REPLY_RSVD_LOW)
`define READ_REPLY_DATA_WIDTH			32
`define READ_REPLY_DATA_LOW				(`READ_REPLY_RSVD_HIGH + 1)
`define READ_REPLY_DATA_HIGH			(`READ_REPLY_DATA_LOW + `READ_REPLY_DATA_WIDTH - 1)
`define READ_REPLY_DATA_FIELD			(`READ_REPLY_DATA_HIGH):(`READ_REPLY_DATA_LOW)

`define HAAR_ENABLE0_FLAG				6'b000001
`define HAAR_ENABLE1_FLAG				6'b000010
`define HAAR_ENABLE2_FLAG				6'b000100
`define HAAR_ENABLE3_FLAG				6'b001000
`define HAAR_ENABLE4_FLAG				6'b010000
`define HAAR_ENABLE5_FLAG				6'b100000

`define WRITE_REQ_DATA_WIDTH			32
`define WRITE_REQ_DATA_LOW				(`ADDRESS_HIGH + 1)
`define WRITE_REQ_DATA_HIGH				(`WRITE_REQ_DATA_LOW + `WRITE_REQ_DATA_WIDTH - 1)
`define WRITE_REQ_DATA_FIELD			(`WRITE_REQ_DATA_HIGH):(`WRITE_REQ_DATA_LOW)

`define PACKET_HEADER_WIDTH				(`SRC_DST_PE_WIDTH + `SRC_ADDRESS_WIDTH + `DST_ADDRESS_WIDTH + `TAG_WIDTH + `TYPE_WIDTH)
`define PACKET_HEADER_LOW				0
`define PACKET_HEADER_HIGH				(`PACKET_HEADER_LOW + `PACKET_HEADER_WIDTH - 1)
`define PACKET_HEADER_FIELD				(`PACKET_HEADER_HIGH):(`PACKET_HEADER_LOW)

`define PACKET_PAYLOAD_WIDTH			(`PACKET_WIDTH-`PACKET_HEADER_WIDTH)
`define PACKET_PAYLOAD_LOW				(`PACKET_HEADER_HIGH + 1)
`define PACKET_PAYLOAD_HIGH				(`PACKET_PAYLOAD_LOW + `PACKET_PAYLOAD_WIDTH - 1)
`define PACKET_PAYLOAD_FIELD			(`PACKET_PAYLOAD_HIGH):(`PACKET_PAYLOAD_LOW)

`define READ_REQ						2'b00
`define READ_REPLY						2'b01
`define WRITE_REQ						2'b10
`define MESSAGE							2'b11

`define PE0								2'b00
`define PE1								2'b01
`define PE2								2'b10
`define PE3								2'b11

`define PORT_TYPE_PE0 					{1'b0,`PE0}
`define PORT_TYPE_PE1 					{1'b0,`PE1}
`define PORT_TYPE_PE2 					{1'b0,`PE2}
`define PORT_TYPE_PE3 					{1'b0,`PE3}
`define PORT_TYPE_EAST 					3'd4
`define PORT_TYPE_WEST 					3'd5
`define PORT_TYPE_NORTH 				3'd6
`define PORT_TYPE_SOUTH 				3'd7

`define	ROUTE_VECTOR_PE0				(8'b1 << `PORT_TYPE_PE0)
`define	ROUTE_VECTOR_PE1				(8'b1 << `PORT_TYPE_PE1)
`define	ROUTE_VECTOR_PE2				(8'b1 << `PORT_TYPE_PE2)
`define	ROUTE_VECTOR_PE3				(8'b1 << `PORT_TYPE_PE3)
`define	ROUTE_VECTOR_EAST 				(8'b1 << `PORT_TYPE_EAST)
`define	ROUTE_VECTOR_WEST 				(8'b1 << `PORT_TYPE_WEST)
`define	ROUTE_VECTOR_NORTH 				(8'b1 << `PORT_TYPE_NORTH)
`define	ROUTE_VECTOR_SOUTH 				(8'b1 << `PORT_TYPE_SOUTH)

`endif