library verilog;
use verilog.vl_types.all;
entity xilinx_true_dual_port_no_change_ram_v_unit is
end xilinx_true_dual_port_no_change_ram_v_unit;
