`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EAEQGCZzYROHaEfOaLnvBL1I+CZS0Ju4XSUmHu7loEDqp76h0uZ1eZhl6pjhKwUz
lKpkmajeVYURzjNAnc3+jEzhXca0yuzl9TwbO0kvasFme6t6dzvB6D+8y03AlNOV
8piyhNnKRU4csxPgkrJG4tgS/RjiyljJaqklHvSCj/kdCRq1SR0gP/lAJ+k9K6AX
UNtZQHrB8aMDmR5NyV1fgnUy2i8b/S/RW2lBL+iBwjoZIsypby3gUzU2tP9KITmk
//bzEseUdaU+I474BrEnHq6R9SaAzbHmjZq6HyzmuSHm74Yu3B4Fp296QwYruVXg
pyUN8YqcrNmT8a8+yjlsShjdq8yJt4arV8XwSO2N1x7q4tbDTeYXXtskCHlqfYmH
6jodu8p882bXzMznXDEltYOHRN4wBWa5qfHxSNiIrmcZ1ih9Emoz4Y5WGwxqKSW+
zzjG0iai9RomcTlKSviGPULb2mLhVhdIHhSuIdXFrO/yXJryLH6/+mh8cgBg3NOq
S52nFUc/yVCTZq23XGlj/DayHRxOgJMx7059lNtFixQFcTxOWg4a3zS83jFcO2Dx
FhDHKdl/JOiUQLV8rgE7dD86rwcticv+F/KDTbfla+F+EsVpRbbhEL7gjF4I4rEF
1GbmC93qAr0Brn95/X5TtJekoYSNejZAB/KUgxvBCKD1pEp7vwt1+eSBdhFjtlr2
WpjS0kcsLwF2w1NvzJY0HUsh1jMQon/5iNuutBQxRHT8mIYK/lGKtyIoNVZ0lQFS
gOCOZKTxe5qp7RCiLIvfRWZ4QlhZI9jQp/oPufCd3zlnCfqLzzNFJy4z/EVS+pWO
CJ4osen2iacLhYDE95Yac+W/Q+f6BzIeMaNJ7xKKn8K04Dad1FIKcDIIRodICh+w
SjaNiofvNz5wSItE7+THvvxTc0sjdXgf2GTzfYr4JOmzPw2itYxQ9KJR+O7M+bu1
G2oTURoF8C8MD2e+PUlhqwX6STvAN2sr2LNtOViGb7uPxgxeETyJFjrg6DZ3UgkM
DrYg8oO1LnGAyHTqDlADCCy1xXqPnquFh4hEumoMiZ1EECKsayBDK+SaVn+MGUFE
mldmMAGl8azfMmHsNHZFGhDwe7uuFiGxB5CGm2srs29N3Pm76A5OrNaKOzPdD4LB
5ojBFQsI66Fr1+5cCcA7WLDRL1n1yZqyMBqXMkj/+zegZI1Ovdkkq5VpO041yOZG
Yj5+Iq561nsUhFE67POsssrXrJot5I4Bl/lW+L+Pc+e4RaJZy5dCkBvk235Or8wK
EZoK7Y5KZa8A/Yof20ZzWLwPrDlj85zkqJiCfTRpyfC1hgDiOiGlzjwHefLP4gBP
IX+pakxlTemM70xqe0eyVG/XVHcUIBJy9/pDRTnlGjvzop9J30a/ZZYxL/m+9sec
5tb7UnayISPGksJJ+DxvBAq4bxclE5ZOaRPmFiYZPqZt5QJDw8LqcIQIrgnlYUkc
aPkyztbG231ShmXVtxUB0J5TdJw2OhGea6w90QyrxEjnwrkV5gkYKc9MFWl54/8o
55inicRy8jQbQ+1ehIBnN521+urfBut5mlHz0L83kZhY0pve5d0R9u/r6gaEHf8g
SdMbs2OFTnAkYp5FFPcrqsvH0iprQuCFG9EinjnCCS2lTp48VGf2b+qAJS+XY5MQ
mZV6Yx7i0CskocqJpA69jefq0wTP8FaR+7WI8pXq6Pywa6G2LZOYcW2l00UqRZsU
HH57Nrc5aE7pszj8qGNWdJFMl2Eb1Lu0JMijGh8NmIC/9jCxH7i6oml+x/Ui8PET
fA5baPJwjgQx0scORbnyrc6SBTjGewAjzdXFLO8nA8zQvZiPh9rLz3UD62Fh5QAO
o1E51k76WSHEYj3PfD7G3NrBtF0Qr4VIL4R8Gdezoo5sFDWxtBv9TTbXJMAc1Dk4
+WbTsjFUuaryEbLeV77i98js+9kTaaOBbM6gAskZFWGkNMj7p4jSHukO5KDp/ntu
CqgMwWhuMsXXsr1zCd7NAtSw+OqoJ5LBrK+gZmJtRH5Zs+Oi2+IlRUhcIO6kAQwv
yya1C0eZeUNBgiA13K78nU3Ub4jH+OZqlxy0MfRIYUb1lNzO0Hgh4Qxt0mrlihL7
mN/ZiYBxALFv0FN+LK6qXJT2lO+kT8+UElaP3U1uaCvaf/29mIJLZ+Xs0YS0Ub2q
zEnYGxC77UwIOnUsbr28i6ERdqfv3ZEr9az0kbcR3Ieb7xoQNoXTGDgc5F9JdXGM
6nfzTB4LgKpuJD7OhWowYiTFY/Qk03AAuX+yzHWmk4fC7HmRB9O6m17b3xx/rZVH
/9nSzelZTSE4eZWenxeLL9cVuf+7MGSmxgIor7wyXicyNwR+YtqhnypMYFXdjAdl
g4nrD9B90GMr73v+XHoZiceyFUHLX0S1f1uvBI/Uv5iueyomeMSYlfNOqRzEAJzo
mUijReiYirrwQFynqzDTjvc3URbvpIWEwigGYrKtRuHD8aCu1cI5B6gdBMRfjI97
8ALemtYrRDirwxlfYQZFqcp/mVX3z4PAHvyl6usfcm4FSudbd1lmldSKI7v8KGzv
PV5j0eQY5SlZuCfvydjWh4G8/Pc1BJRzAJZsPFS16WwK5yVzj1f7MzO5SjimoiJZ
Dw5uDZmlnbJUA5K+ALTokai4BrSjTUGWFbp/P8DJkI579Uuo27Pg5bh+DUcE04E2
X2dEK8KMqExcrOb/VtHB2dYVz9jS5N3TKnJzrXFdlfJXJ6ZKIHOnMQaoNNqlFems
Y8sSYpibrdX0MwVRuXF6TbFVg1SyL2sr0UV8rUhR6TkZ5kNVYhv2RoYBWiVEwYwB
/8NIFLk97MreOmk4KWNr8c/zYTEvBSMxDLgad1ZBS3l1HQKPcYYy7Kfwh8lijozh
NGS2yXzqlRPFc7T7BZnQ2nXxMz/fqauNnkSifMZ+MC3AaKI9iq1v20sAeNS/6P9B
Fi+bTb6X1LMZEeKIewPIh87tJ+XP87BYvgammMRY46yXjzzLe2xTLY1cwEUb5uTP
ofIQcbwbyij28bWUh3oLLgn6S2AN9NG3Z75imxaxdac+WCZ9a5/2jQmQIJFTO8uj
nXNhyNw2RByBHAEgYT/BybmmUQHrXLVQVZFoCZJrrFSb2tIOcx0Z28H8XSqlt5JU
IXLT9Y0lI+yZGvecO4vlPdRJ0qrWgjpgJBN00tIs3nc28/7pHqw8GA/4eVAfVH+c
z9vLF5befxxzXlBKVr0gdkGaXlJBU51RBvx7Ji+vsNc0iN1G72UyXRI3JObNfAIA
t3KQIwJRY1+g5mxongr2sFqbDifG9H+hpjSaBB3Mnb3tnko4HCtPbDMf2xmra86V
0eOJ7IG7HT12OcbBAMuJWdvF5rngaMv0DZWus3TBS1hAUZRn7mpHUYdAR8jqev8z
CYRx0m+AdCdaNHLrZn0ZP91luaGOVEY3wkCNhN4TieSxmz8hXEQSI8uifzHlIFrA
ARoHWThhJMs/uMqPvTozeEwZAU63BxMBKYyE34ULBW32eYejvW8syJnZSMInEd9R
ZO+tB4fMhdAiTfIV177/CEMeDjesPQGAOz4i5wvUW88nshhIbF1byq4qcc9H58q5
RO9UEljeGIfJ2Cka/goyug2JejUvWRSt3w3sAALSZvA6TSpJOJ8iEedP3+7qc0qo
JSRRAU0PapBESIcBDUoQdVJaR+vzk9eSOq8KRGRgt9IU/56MPZku+98ReH/zqboM
sMXr149VMQYqwKopP4TwpLEt0OtuPwct3O5WKqvxqiPeh6bmJkbfg95S64KObDEU
wY4HUH3athvr/HDpmCXsmnMgM2lUmxuzQFtNgDO2l0I0VGTg6OR1JeTbnJ+dCgDk
9D6/YpqqpeproOvG9Y24nv6a8g5pgDhRYcW8AS/3cSctUHQiNIeXbs6WRrhDcj/T
fQEVaqTDg5oeJfdmL/Gdg0fRE2Qx0q2KkUDongT1QYtUg1UCD98hc5zQLJBUPWff
V+r04twhAuImT8bnAj1mV8LTiFmbsazn63tQkyEFJqgNdu6WBQKVOvmZbKh58pu0
4lOXcTxS7LCc6K8Ao3h3l2CboyhJJHn8d7l8p3DVBzIqUCNXozxZy27QQl56X8lB
gvz9cX5ROi44ElSYsgRape6Kh0BKR4YqVFCyx6WsmQW1TLr5n6ZMB+m18HvYfdy5
7FizN3lSqlF6EqsFWv4DA/eTNOYIbC428lfzG07IPcOVspTgiJfN2xPHT05vWOt9
eWHok/urhWDJJU9KBJTD7HYT9OnouRaevUga/bA5BxaUQPIKVOugZ9DcLZHDfi6a
A+IWDCve28n2TEL1OJcsCvF496RoWM7pogBFsr5WS+zMZ2uCP+1gNP2s1/uHPEb9
U6zJnZ1tJwh8WumAIUXPHrvBk/oawfC6NCOCPMyMYA+81bQiWbnBh7bWsUFwOxL+
sRM9c/SYEbXtbj0DiEP8WV4R51iSvoctbXAdAhdNT9gpmHtUATRHpgSqFSw6ztyd
qMlY9QHE09SOtaDN8xSP6+FuwhfSKHqppCBmb4+WHYLTw50Tl3U2KTYmA9No2MNS
GBlJfbOOfEzLOaHoutZCuexaZBdRyG9f/R8P/cBpw0iALVdk2DB586XHcNeP6Ga5
K1Yq/MsaCNfR4VY02jLtVT5Z8D7D0X4byaAj0Ax84NwCtJPPZXpxrXdKMejkBHDA
LHDGYyclUf9647PIirleS5PDaPQnvJkUfx8CZ/yNrivJlUux/B2yizg33pQoRg+R
ZEPWqlIxifKsCIvOD23G+LMzQFqqH6stzDKxKUP3aLZIm1Fp83gsju7mXAGq3R/l
DAKlIvJ2LFhN82ExQzrlXhmNyr+KwOpOZPqMZCyECmkBm01P0HvCCT50b8X5UxXk
ZeyeIuek0VNFbK0VCn4yNkKK16EX/UdzYXtmr0kPOGrdXfRkW39c93fE0QqdMrsc
aQ3DwtxQvmOq+fjf4+ZmolOu+3QHtI3UC9EDUut5eFnVRv7Au16ofJb7sLlnTJSV
YDBgMTvCJnFFChNndAY8c3HryvLzDtpJY9VIRuWvW0KCbEIHPxJ9M131axCmZV3p
2mI3pWUp4uu+qcFMaTCtnam/ogequAL44IYgN4nKD+9sYGyh7MhRB/Y5lMFLEfJg
WX3Nd2aqDulGKf0IHytTSxSF2+MgaUd4dvVQ4M0XOTgi/05/0k7Lwlr0Wvg8xU5M
aZB1CBrqzA6je9bXr29we0Ogw8iSP5DqBkvY3LepxLW6NQLYVqO3w1oGw55+gwsp
jmaPT6d1I7IfvXnR7+6cSPgPp5kCkGxKosyOD+I+EBEbSTcldJk9m2GFSGpamMfG
Ro4j0Rzc/UfdkrevhMh6h6996t9AQzQMnUO2oo/yr8JGSLDuBsYUzpayI+RXNG7Z
kUBqFRh5rDYG6IEIx/1gJ6sHlcQFHpSV6wiPQqJ7P9hAYzyJjrpu5sPHbEELPhYP
kNJHTMNjNgw2t6ZomYukTsos7nciB0ObRWZgsy4d0MxDB4qS6DX16d273ZAcVfTr
g+9NyouhenzF7u9aaIFddV5GU2VQbFtYLL9Cg7gcVZoXrli/YQLwb0aemB+NkLRe
hk8qs77vTJBQv/RDdCtnM0tMMOzpDGygzSVNaDNuhLbqjUf6t30rwPXPRus6z1bu
cRT3paFYy7WNimBduhhGjlsFO5j/AQ1/Er+Rjz6kNcTfPdvOHIqS8RgS7+w3LDww
YbZnFpQAa4Oim73KYyu9jbIZ6VyeA1l6HahnlNHbo8dDGtgWImUR9SULE3ZAISxk
pCnGJYKnGdLSh3yVYs/AkVlBmZ/g4zH5h5ZeljPENbf1US0SiRBx3qBTp/QL+hv4
DCYtmAaRKEsPXK8199qBNoJVXVyVSdGh433gWyq+zJz3FFARxa8FvDQ++NON23ld
pIQ8tbSgMqnrDMZj9enu8HklLqNtrfrgnBqyEMDYTCxKFZvMU2woEhNyHBrAMrhr
2ms3zxeP/cfue2htqKJwwd2rEXwKUlqf4r8CPsZB0tJYsb9K6lI+0SUWKzcTFjTI
Xv5Ef+a/jGJf2Pk35B9N0pWyzM0FYB/km79bwAvSRhFvcPI2knn7dGhSiE5PfBFP
YcejxP86dz7lfX/ttP7hQvJV7O1+2keZyNn9Ye9cYmW3DiU801+BNs7yJLKXn6NA
ZUwHTnhdxrHdzIgW/XdkH5ci9ilhTTV4Ug3KhBdaXKDe7oP15GDlP0qDfRj9xgXd
yPJ0i5rSv27/t1vFtdY7c5U8qNhRaWoeKm3kT+Tj/V+ggF2EqdbgiNoAb5ap7a2c
VdMiolDG0PSRHb0tfv/QcbD2dbuMffX8uWBynku1GSqHdEbHD+fkz18PoDEw0mfY
ITB1HuP69yecmm2N+A4Tdru27su+m450uJuOPtC8piky7KrKPyx4KyU8zFRUGAJB
qsRKs02cmgXCMpVF91h02PoXP0B0Fan4S8ecCi9owDaoq6fhkW7JYYMqRl4oV0Zp
PtK2cOIx55XiQdKAwxu9K+rsMxACtGLVjG5eC5zFw9jEfE2J+FxL6CjTAS5eStyk
ZQq/VLy7T2iT+2pQALLG0i/6dxy59qJY6WG0lr+CvdaBKlQc3lGURYUp/6zi/nNJ
QKZ20HCXOvJ15rkWW9G8n7cQjHImUXfgE4z8uRIk/budDL0JQx7PTOamy1YAfn0k
6GyQvrqi7qw4K3aaQ9Y+UyTuGJ9tdJBPmIrBHjmRN8ePhp/NADy5J7/ri+vNgmAb
8O9MdeqaYFWSpPcm4xflJvmamj6PHCpeV/OtC5njkAf0bUwbLaLKTX27bbRuMIIQ
LiIhua9eR3agIYvFqhazxY5typCM1/r5YHYXDFx04mq6ndUJ87Ajy6c7/+YDDgZR
8FHBe3Er4qfMMl7i4Fj3HLQavoazdM+/RmjtPQ1S7489VwdHBNZG8jHAHngW1zB8
y+XM3PHvioj7UTwJtu9fbaaKgLr07RA53A4hWFZiIz60e1kxQpuXY8YMycijBo9f
A70SOXgi3BS7T0293QnV7LsxTRmGAGTNuRDznmxIuPJVSglBVVkCpIOOM8oCPRaf
t2RqAPR+wce2VNPQUtltzF0+WEJ8sljxApITw1Ps87kKr8gFiDWPnjc3lYrfL45j
nXm/Xmk9rYaz7ZFz2zphSMxLllq0yISn+JMSN/pv8C9AyUWWPf0K21VIDzaF0ixz
lUA2NouZFC5eEj7uF8DBJ6ZdCrQnh27GymjzxyI0tjEc8SlXnrri+y5gbiF0UTWZ
gVSP++UMRYRMUS/QO0t570sWoTuxRWqJdqTF19lgj3Br2VA7pSnUpJKCW1owdAOJ
3A596yfSo5e8vLlmo/og1GGDmN7NwivgK+H656pqT0Y6zQ8W6q9U3t5YKvd2+LoX
vKiSX0+fAfdnaYCP9DTbJQqH+roktiS2GUkNbTi/kYljO2ZQQ/MGi7d5O0hqeV0S
oXybPP/I1ieZay+AFjGBU+pzv5X4LswW/euWTJiMkyzhUZfdgH9kDPgwIkFyBsHj
T7JfkFakXNCkoZjIGGAyxw1akwV/8jpAvtFEeIlzLsA6kap6JpU860hbEs22UVWZ
9IAKZQPYQoOgtnqj1IGvihQaaBfIaffnrORj6tpdSMaO0PCofeeI+8fQTxE6ne9B
Drvlc/8ERNqPHQB/YlgyWHP5p0gVNWwmE3i3BKI30txn4Ut2YSuz9bVp9b8pM4ll
d3uO3gyraR+pPMss1S2kh9TcnrUjSGWbB0FjJc/io1N8vYgz1mjozn3GU8Pe4kUs
jK+mQtOgdmfQMoAdVDYaiyx+VSQS0WrtlH2jkuRt3qMK740mg6482Bee1isTx6Hc
t33w8Ba0VRs2B33Iw6IYG7vD5zYnn/VtlPYhdmLHB6PMM+9OfXoertOG9yjIAgd+
YRZwC2rGoK8kBn7lfn2wonGpbymQClutrAuWTRxB2L9IlLjLdgR9BsKqjrYfBvM/
4uJ02gQkU4af4XEDx+UPu4t+nKNfh0axs4Ony8GIywPpVmxwHvc7vRiL8HvHiCoC
9YrZ7oczqPoe5fuDH0KjkPM2mtEqyY5t6O28LJDfvz2+7fU22H50Pk2vE2k3c3fT
YcU2xVZqamBQ4Oq+pOlpJN81tf9HIdOWPNU1CgSCkkBNdZ44EAya3j7W+kj7WP3R
pH/VZ468X69Tw9PQQskV45eq+NnjpIM2psxr5EEOwDnM+fJ2T1zb6afzLIx1jkFL
8bspTp5UcgVEBQoziVHNu/UEMMp8PSPOtQ2kYzftchA5KHt9478EMKbCSFq9nCOn
1CJYd226WtlIOOFRR5pt6Ha1wV+tIIXsEC95V8OiDDpc07xh1hjM96JyTkCMiGjs
R1CHHpGw5d+2GAHz1bxKHaz3NbW2tINaLCuSAnVX25zZijBXT+CRkP4SlSEbBW7A
LLrlz2gx+ildoW/+Ew9fMudVNDEHUnopMUTKnA6NGMRl3VFyoSKQASGuZaELZcyo
a3CkitQrL7XTcbvNBL1l7hV1UWVCepczPqILAMdeTvFxhaqM7gFovnJ2/zshEsaJ
n3AeFmYFg7pUVJw2RNvotr+zR2OdQgjnBNFI6hDeAHAKX6mYcMuN826BiY71G6Kt
Qg8TsNwXB4MkVwMHM9XhzvslrUZ9ROAvxD9H4HTiADUb4ROeISClwBAhmG0FQcxf
ttYh0MOfzYbPlgE8QM4h48MlVm0qOZDueeIqrfujwHffbXfOjiHKrd1+3lMR7A+u
a9JETvYYK6GEmyNknDz/RDi4SmxgYjbsIq3W2U5zKcm4Gd72HB4X8c2nV5Cj3Py9
1jq8utWWW6CyXhWU0o/ao7xwN/GGOE0gWU7cw5l/Hwxc1bC8ReyenxCwB2VPY8Wa
iUqUOkgHW2+aMGz2A4I3us0VveVYMxCYnsp9DnXF11/1axPerljWG06yQ89X2NpR
hWY2NocIpyCYJF+yW5DduDCiwlQVjrvRPeqZEZKljfSRhnE+CpCbv+d655gbydd1
L1vdVeKQtbdZCKaJHQlkYJj5f9cm+edawIzWNyELCUw21zvAnhTcu1Jefa4MUhs8
nt+wWnzjKR5TI1apR1VrKipOMcChBHTPQAChuO8eQ/DjTJ45Te87geU72ktwsmei
/q/AYsrqckVdmLVFZA3bOLnFwzEnoW1+pKJO2BDvQfXsypvP0kDPTf5UXOGwh2jJ
Q6/4xEmQI2oqOMCSyr6ScVSpGtR2a+COzE3xFjYb6HM1nreS9x7r6Mv8OBbur92Z
mYgt/dY5t11qeqm84EeGeyTP6BgHMgzK/vLa+2fVoP1VYSZ9bE4rQXS48DPtab8I
f3JIFNGJ5GVf7PKfRqoTS8Rx5lpwf8/rOk6Rv3VwIEuFNDAi0kjg4giVzA573MfC
7XPpYVGGuOSUfOEStg5MtfrsBChHJRG+unYccmH29pTm0fvtvXCs+fm9g0bqoGMw
mpW6UUcGAE/9k9iVmgRHgv3L9jlvpFLKXr9T/eAdMU96r9tiiU6lOVZTc3e0037v
zy/ssdBsLw/rHhEtDNDkqx1/wCf2VEj1+Vf/89/TPkqcaUWOd3JpjjQZLOGKh/8e
sfq/rCKPsfqypZFPZCV/OuTc2hXj1x+p8s2dDrd/6xE3PQmt3/X1pt9LtjOwFmGe
MtXTqJiS4enVLj5PmXXnYj0IeJJVNhN/ddAFkOqtD1L6Rh0lalpbeHkFY4M8D8IC
EGjE6pHA/cYr6DdBkCKzgNxF2dZkGuXUbnrWTM9y0+U9WmsWpDSbJMv/W9LE6GF3
xP9vUEtiaSVnPw2Mh9v6bXRoKiuK9mxjEsIEOQzxPdiDzkCxAGkuWohuv2itmolx
pJb8gnEZZdWJCdSfk89zB8wu6ZU8wcLLWBqZoOkZADA6P4ZriQiRy8Fg6X27Qy/Z
f4onry0fYpfig7Rq1gAe7B/PSFw4Z9KIret5JFyLi7o7KEVsgtdWLgOWe31jz3ae
hW1e4cSGOjy4OyWoktp7IqawxkfIlUWNTfNWR3yfkluiaBZP278W+ZqeOZgq7e/0
Q79BPrMHMsbbl9g3Ocf9AXSZIMdpveAbP89i9LG53cuEB5QhjZUrg6vixfgL+5Mp
r0vM6Jv5B4uu8JopauyYvMBZQ8PN3ISnG2aK+c2Ec9X94CFl8f4VDk2oLkxt38LA
F1lgolalhmJ7Mla+GVfXUunXOVJv1gG/6Uc63+f9gVq/9LIvfKH23EIjocBtdTgQ
DGVEcDLIAtQ5kDutt07fYFKz8b85tmaTufy+0St8ISOFcp8kpW2xrB3M8OICeUuo
f8HjC9pNWU6eh2NkAD5Yq2gyyh8E5p8eFpQaTHsc21NHtRdUT03v1aLYiBP/R5oO
fkPvcDaJkpQRKMWKDZfWVDf+v8hobFhBXbwsYZrKe4b1Tw82WYRHTwTEKcvGrAlv
+sMSkJSQy13VeSFb5rWPrq/6aRpoePj8AsffBKp7foHMKsc7Z2ueFAQg20yXIYKq
Sckz30S3oPGM8FLOvX9v4EMcXwkAyK5aplmIbAxGQqs1CXJTdwJ1PW+N1RXaZcgp
hU6/fa+7v+FhTGMEA9BlShgVke/AN+Tqv41DfjZP1biSrKO2osXzPyMto/04G7dj
aWot2LrDAN5GDD1JJAD3N+6euyNrSEdFwlNirRnNzcpcF49WBz28PuL8Tj2MWxRE
SzbKuuSIuAaEySLEOceva18+rsEZgvzM0JKc7iSWrIVhyjBMr1ef0xiyXRCrUX4Y
1ekgfNXFhFN9sjDvigywifiu2sZJoLYRP1ZUWju1krgKZ782z+vmPLOp3tupxK6j
EA2WjyzKty/4v65cUQwCa41bzBaXjqSwsOD0mgqMTHMCeB0Fs6JmfRfraG1agXCN
T85kn7ovYHkl+SBNdPRvjGFYpuPZ5xwrj9QoLhPq3CEtSWp7utX1GiG3C92+DRZl
Ez/UdrfJpPPBJHndKED/Pny2qqPfz0x8fNkj7DS/sRuR0aeSunU9HArRigagE3CS
FW+QFiq0k9XPsmrjCRnsttQfZfQgRJ1Wbkx9EgPx+o51knooRt3loFdd7NhSbrdj
PxQ5IuRtkOrGVAuHUvafUlSzxroQ/2pYGIR8YP3xQFuyL1PQoj8KwWOi+/L3EyLh
HTpfUUKrb2mNXxTjgOkWOoxLOmj8qkkEWWZiFCkYObQhKMUW1fnUmPb7aEssp4N8
4XTYVpAii7Xk6brslaSgqofa5GRtA6xEFpAAoilKqQ+03tCLs0eZnn3C1Zgso6ck
TxwysyP9+Cy73+6stjmv0D9ZcXsAngbXl1tgSnBnIwnCAYdmUGxPeZiF73gmbLLq
SEs1LPff3nlJDtz42D5hw6cKbJh5FSq38n7V0KlKRo5sYyIUXUDkQ/xJ6y4xa493
xdPoC0Qc/1bIWrc9qGIAoqi7pYi12nHq4eWtH/QhMZRM29F+KH9ArXIq5GTdZFjc
g3e5YKkne5oC4tlvS+8zYn0m2ScCVRz3msBpSCmmPYJj7sUv30+UsUsQOPUcRUlV
czsBtJpblKftBgB2BNDUtHTbgznnTG3BaGFiHyEUlASUr1A+/t9UvH1SnkraqLlY
nfbkp9p64JqjSPe6+NuU2of55R8erGbTkSA+MKxFlMBmdUGoVGh9947gtd7EtcZT
mz0z1PUxNCZ9fQoZi3M1BIQOVYWUptlmJv5Qux6W81N6NoMu0mvf4Hhh46TqpRuT
FHz+RgbYVQLXkSFVr/aHo92G5inBljzhKhmgw5rHlOoTO7sWelno+Ul8PnELlGIb
vYIeTSgg5zWO3XoFBleRH4yeBKvuAe4HDbekb3M+M1v3uJdJipf0e6VFXus7Bb5x
ywAH4KcsKOZrzkJvdZu7yC9Ahsmj3J+WIQAm/yaBMM+pVMHZ/XZQaQ4HidOfOqaa
LTqOIKqbtOB/D3LxtVBR/m8ppNkHxdp3k8/DaGnV2qw6f5Y87HsdeVUAJ+3mBALB
/vrSSsR2Aqs1ZsDmIColRHr/QNdXjpMFbueO7D41cLrmLbCcNqDU35wd2CwJ7dEd
wgIZzCEUOR03Z20I1YMPcnCFX2jhkPVYtjPyfvmlyqOlAGZBL5Z2/+4JW9gn986C
Z8YSgTM2injXHNrxAD3Lwk+VOP+XWRLPnLu3T6wwKrS5vNJldvpZKnZxvSZj8Vec
O0b3Ri88RHPyjotDEetnMF8hCr16JMB1I9RmPndpiZYpv9a2pwYMZ8XXM30ltwrg
7FjS0UisJdEUtew0kb+WTRmnwTYngEnJcaUtWAXAcjm+KPoofSswThtq3YcAqAb9
WmMqx2BbYU8it9JC0RRB6qrms12qyiZJ9ScKsGnh7ciZFzc385yH6wRRcHbAqVCm
/rXUBMQQCicWuifAF34FrKG1pC7+XmT4LOAdFG3k4vPkZOO0j/4eqx/ZI3T2Y6fk
SVRwrWDToZ52Zx4PDIUXruNmQah1Sj5ShTq05fygquF650Lm5QZlMEdOUjURHvSC
aUpOBHFmZixjL8je9GOyMd8jnpJCaXf8paRoPBZqFnob1v8n6Ow4VQgs7XjcRScS
vOreQv8VvunRvc3yuqiQCqqOVAxu7jC6A28qP9E9Lh0Uobldin8hY48z4pSLwO1Z
I6pn2Dz1Ej3UuUKJN0ZLE30W2Ae7MSbFdKMba0J/20Yzxx7RKm8WOXyFsLOKQ0zN
eZu3ESKQv08GtB3/UX6X5Ebuuy5k3ooaUw4DsWE42fMlTi1+qHqArRxUTZh3mcZP
1ySkNIC3CYzVgK+ifHRLmZ72H4IydqLvbVuKzElF+JKYZlMYJO6s37gSGCtIDUuM
B+SCJz+u9HQuUpqGXeEUzhFVk6zxcmVu9aqyybPbMMZ+dn0IfPRblNRQGFTPXUgN
WbwQZszGM5WvfZwVrCu7zPZUyNh8n71u+M7fO6pIcPd2S4I9OsyK/9Ez7Me4A7cV
FrCCMr+czIgGAdX4RW0dS8f5YGuxGokZUNDt9O7gnBn4YzJZcGjhXqirKNEt3T54
Xskx31qCnRZVzpJMj1Pa9O8Efgc7gHqbFppO604i6XySatLjqor4KI4gyAVonPl8
GTvz5eftvrz7IktHF7lzDBrLnz6RfzSUNzW3yYtSxrwMRJMfAhtawcKN4sP8w1Dz
Wu37Ey5NgodNmVXciE6MMiYyVUyBn10eNXGepHAm17yKYcD46ST9RvKtjqYM/NmS
isAq6APEo39aJfD4oheqJlx4mCFwk6DYklAs1BLl54pYTEWi77N0Y/HYgRhxlwME
O7a6gy2ZvWgBQtelW2cgnwlrtm1YLGS7Is1DB7sBHoANWAEAsBCl3rIwotPzvshW
25obLQyutRWscPHAjfLE8x1M/deHLDNWjpBYECYgT0WzjZvjgmMqfLpCd9RaQklf
EP/9kvpbuxrkrOuZ1WtTih/LM49iYmZoe55jMe3labMLHbncp8lsxHalrnvDluxx
8NkeFDm/PdtPlGaDjPxKZqWQ1JBo++EU6MJn3cEh2js4b2kWebPRSb+AIoqSQgsh
X3FC/88F5CAzJN5tLBTff8sqWCWvPcLx5SQwNW83m6nZ9oz7No4SPUyi1Apsztmw
CWzL2lGRqy8rUrn8q8caajUptZWbAb3qDLQ0r44ndNCw/aIEfc7XFIHcIZ3oZTF4
PKb28zLoOL7mN9MYTrBsihd+NAsg4NcCb97Ntdv0udHOdxGX4sn4JH4/Jz03jj+w
W/chV8AF9gRfHD/FFCLIEbq9OA4sLkqs82IAYcDR5Pu9BiUV9nW21/6LSsfAkJCV
dwJv/32/GXREWiehiIeoGuGLq1+5PRldwx7GvMu+sNHnpyrZNuR2QDpwak7uKZzm
64bHFvVjrF9Xw94+hb7my7W140rOFtokxv8lVMJTgArVoz8GiBAsILxb4a16q7AN
xAn8F19YSxuyYHhSjahEULsnLxWLvQ8+c2eIH9wCzX2HHfJ7oKhzIjRuHNuXddsb
G4awTHGCEK60zZFdZpOgxh1gpQPOoM61UhZ7N3PhGE9tt3i47p9/Py163D66uU1A
RdQgg6ZME7hNi4HDyBhYOyDZAWldNrpGCtluZlheKhv6jsC26sYHLeOrcNs6/xdk
OkrGHD95Lo7eGvSinWRcd5zd1MwnshFjO6Mi6XNcaWfrbIjFoxN0U/TrAmse0rph
0SyXXwqB8COoja2BgEhbAdJEZgx+hAgL4zL0VtUfOL6mgtFCcwWvlbcvekNfgs+1
WnrIMw2ggufeeGYMFyJhcyX2teOH5sQjWpiuXSX0omEMB29M+62My5iN7K4xCVM/
ZUZpHddRaxCj5MqgqInjyea/2gqY/Csgem6UqY4zIa8jeDeafjsIPTLH0TV5R4q6
1363aAcN+jW7+1hCY8loJu21R+OgbRSsSw64dhScuq1TOD//8KTRUzSOvqJh9DuZ
nb+pbM8NLJeXMVQvokzfLpjBbn4US4/t89eaE65k8YOAnbFMGzD8Wq3B99A8lhnK
Y/N7WU0TeHEXuqBH6YmHc07N+udIINZ9ddouPy9+rY0FwjuPTW+suRuccUgI/v9p
sBCHCP3KjQIFafGiHstcYOsG7mPqIL03W1k/tfkHcrNgwO0jDv4eQ/8v6HWLuwGI
K/r+cuNZtZihcMJBoAoh1pw2FkAV6Q3SDzAO2oUnBtRvgkkRFcmI08SW7yFyRuwR
niGl86l43NcYLukforGfHTXSy97VqgQNqX2L06XM7JyeVyFwh3uxevHuTzlA+sdq
XYBYDVCB5hu3pIs1Z+pzZfulltC3CZhYVwH8t4fMRzZppsr6uuif+ykOAyz7Dyo+
e+z17BPr0pQ+G7OGbi0m89T2CBEsBH5dXmg4uqUeoT1+b6N094TWDWQ9BTD7oDr4
q8DDbbiYtstZgftwEcEVWm0QLu55dJLbMADe6WGR5t4UzpEIeIrBrzq+weonMeIl
JHADeFaOUISK0x+1Y4bxf0Rqotquhxmz3FUNcsi7uW7uI6wMBUB1ByY/jjxSR1gK
aA0G3u57iDcW1sp1SZJ4mRF0Lbeke3po8LEy1MIE1SQpX18vlVVyMBYrP1FDqrlS
F447/NS42mRRlay+ERodbngm7cn75DJQokXzW26tx8DRe5us7P1/okw5I7HPvMD9
x9xyXaQEiyYAgZBZ2L43Y4QcALXdqnUC16pHPmPG/Oxl1MmzpIyocbCT3oHGnJ8n
eDtERHx8ulSz9tQRoloRAwbT9d0AjWYzKUh10dGy5Bd25V2FDzDwyasjqjxuXFeg
XdqRT2A6pQ390FzzNT96k2dSHE/2W/5v2vXSe8btKUxPpxeNAAs/rOvwgElLz2b+
eb85ONB0WgM/tc6YK0vVqh3Ilwzcap7/0XSgatUFtPWvteV18N5hR74RBg7ab74h
qtcI3edjrwARw7pt8NdhH+TSW1zs72g12QYzMlNt8PQBghx4DTdZ17Mkiqz6hrB/
Cjfb1hIznxX9u/sbU01MA3WsPjWvtz8SfOrrqS8+hxmxR2te0kkUOvLYcUPJJW0o
9YfU/npGxalmAEZzk1cymJRWSUxyP/fYEzrnebtE+AU0UwCuje4Pe3hGmOWVYLrW
lATyokojH9rMFUZO69Pqwhc0rLrXia482j0W9HAy7RfuVipu0fxEeenmLMi3+0zV
ncaGnebxGZ9lS5e1/C9CAPbg01dPRoHI9TFpkSEBm6BFhIy9JwFSbfUxiVHSNGEb
pjydTs3iap+8S0ZDpFq+CjNatK0GAhiTtJ6DhfCWfiPytnhD4SJXUN1SBcQTtzak
6MzdKQpZ2thzqyv2sZOQwhSd5v3A35Dq09SGJ3ejVhXwXHlrW1HYWiu3zxzwNiaD
czjyrh+Ezgf4XChqvfNknI3wjq80GPG9u+oJYJMXRxbZUxt64K4v/FrNROukIsLO
Zj/wETpSe5qAXJgj1Zfpektdn4DB1XKzYttmCcYyMrp4fHcW4vBVHnxwoPlKApQQ
Q3POpXxhaFOCkRcXmD1+DgfMNHEuxMa3ubi3D9Ilp6QR6UpMy5jiZeipHWoKC/My
Ar+trIGEwRRVQqWZkLtkBnqW+NhnNrx47w222btu73kcpW9dQ+tJyIFG2rCwoL/i
NRyeLrF81k2e1rS0k8eDW8rO0ZdZx9n/GgvtdvT45Bl2/RstdRIw6rAg+gyhZH5W
OjC7db2APFtgPg3KT8H3SnaijOspR1Vz7/OQKwVkqhoOqpEAhRHhYp6+A/VmEgtg
oO6uBv2sErVHXQViAU/uRoi5W8Zj4SPDZ/M73/z0N0QUxP2whWYS4RUH1pebdbEp
IfOFNgHa76fQJyHaFHPpoMVpxLDoaSnZ4o4m2fE+WFheXhfTE1XhWQXCsQkN0yMi
76ZZcqhQxqPtCuUbaybhvFaIof1vpS01sXB7Qol/lSrxQGfq6L6qUiizPQs9jDRc
6Kzd7OgBrn4j7EVGoMr0mm7fbOKsnh6Gim7eBXaDiLeQA+T6dikDu7b1aCAD1sQG
0GvwzDIt5dv2EJgq8iVour6UsrqMyTZlxf6+9F0Q4jSVlzq/H4eAQfFirfL9AuQj
KbMR2XHFWdJtdPkmguTV3oKSGHl1eg34KJN8w4tEwQ8L3PrajpDagGLegVGMkm7o
ynfHrOeJcJpaZXN2+OPTSPR4JSobjLD6kz/EIaUygkZckuBFwxgG2wElZrNfL0N9
3n4i1iAz61o/IAKJ10/ZTt/yaYORkEAQRJ7bGmU99MZK2cL/4JK+dlGN4TxiaFDl
bauAcswe4GJPE0EXhlRVcuWns/Wz1bKXh5CVj5kxXOxHE42aTz0APzROOWXEcEUn
4MaOLQdApE5xInev0nmIw1NLVCFUlIiylG+vsvvcqBwYbaX59lTrLCTD3+tb1CSR
B1EA2C1wPE/3rIv9y3hiFzkZXTN0Ct0U7oP4hC9mBx6ipyVtKgiJWe/jRmijsT5x
V11plokHwoYcyKD13qaG2wYK4nJh4BUyXXzMehj3wSzQBlXxS9zbObC9Ym6/Z+RM
tomLx4/MZR/FZqh30Z+/BuCV+oMRk7hedzEYJIODSx86jYPNhXdPcHkpIvIPvTzL
BpEGKy2pIoyYRGDdn/QgtPt43rxFoi5R0xgxOyk8/HCev9n6s35SwBNyr178UYxK
FAyXaDBOrusi4rDnaFHm+RC+qDEU6YRoLXV/wjnfS++LnfyxPmOHL4bieAuc4AUN
kqA/HuzyiIbyJY12o7yl1TEiSd2tbasZt+Tp2kx5pYNQ1Ce1ETMzQlBcL52FxnL/
og8Fd5uyQoGjSs7xLQxuODTP3Ry2KirXuW1L+rs+sEC6EfJ0u8Pyg5pwNi9PjZZR
FKsH9wUZ1ojT0ZPrCJ8jMEdGFiluh4dhFhO4BRDYON+X6j/AECxTJzULxTF9fLIN
tvZHhBwv+2Zj++mbvsjs6PPAJJKF8ZWsJKasAt4TO6SBo6H4kU6d0UOuBp/sKtux
DvGYQE8XzMaAH5xUxJV72KhBqwyPkl6/PXUrHSzf+Ocdv2+j/P+kZmCz2TLztw0Y
GTykIZvrLDXASJBvSc0wF5F2pj1b62HPbGZKHsZuKuwjbWWOzBF5PcKQSNBP9z0H
xX9qbyKBdY9t5MJzpI0+TALb8SB/d9ZZbOSy+KRu/VNvCBxXF0uHi/yHAHqHQ+5L
dM5Wiw8BveYtwWBHkBNQlDdyBLkZRjRHJcFr8l9aPEaG6ajSYbMrXDDjFiSQ9pn6
0RSgCmGCuDMtzomo+8kEfmiBeWtIVtfGkvlow9ST7FnBWLIAIGWEF2m7NwXXo0+Q
o8V+P2WMiUsP0wcvRat0XF+B1w6y5AK+CT5J/o23D2Q6njefk2yzJPKDCNtdFZ2d
KTs7roulyQr8ibYDM6t00ZSoM4olnFn/hCAaNx72zcxlMdOU4WijtEO8eo2n9aY9
Lv0IeGxY52J+n9NisU0wjKeAZXunnPxUN4VDzvTC+Bt61hBUkjz8kz9Y28dTgKQ6
QjiluTcpl0uXwYtWTdMSDmNVLO3NSXEIbeppJ1eees1x+jQpZMKr8t3vrPJ8FbTF
trxxWcE81EXqmtFf4HBPvl2tcA9LYigqLfGSyp984+R/5n4W5rOVSrzspmfF/+Yf
Y03GQtFd6QaQTrynjmIlPRrFTANIGHYIjaU06WYeZt/nlfKK72czmLBPCoMBvjjB
qN/CMudQnqCoS3xsOOlQoX9/aGGAUXlif6Mb+UX0rlr0qw4xPpjaKe/f68yYveJ5
4BqV3k6EdO0tCmte7KyM9DcO1gnJpz01ow9eP8PdJvClU/LY7QXtH0kOXlFRBs87
zRM1IS6xjUxsZF2KpSQ1Nla4m+KiM6ppZQim1VXJNbFL2IeIiSTC0fBsC6fHwaL3
C+NPjvfXUgmN2vrQ27r6d+XXrQ/6WC6LlUl0EHc4p+OFQpGD4yXZfOYm2u+7DAyP
kpIdl0osUho1v872dyGrxqa4ARq7bTTO3mKtVtBbaKCgLkpN8dqVzkeCDhX0trJH
La8cKryij6VV4uY2LtXoWGWMB9WpdulqCiDCbVwJqFzUUlnV0aHuqUvSmxgb1IP1
F6UtbPvG1ATg7wqZ0gFfl9ZZvH/M4wno3aPTfvC+DzIAXD+c2xGt7T8bh08n2UZx
hp02lN84lxclQmAKxJAHEtFbzcYOHIQ5FijTjlUr32dkFxpYDNQnXhIkW1P2EFw4
Lm3YY5OTqW8Ax9fi5fWPfLpKhMzO91FCtaG0jsmhPQe0wP0byAF6YKO4SfQvVzAM
kIqd+WoCj4CxcZ2FImGQmX1SJC199CD0fSOba7Su4NKAE8uB//RvAKm/8h5CEI/Q
pwCI5EXm9Ob3h9rtTHbMtr8JkxjFTEQZNfMbuIvztgCzOtOJQrAKYWFUn5m65jHj
5HkstCoYA/E4J51f5ooMLYuGliMtxHpy0mndZcjFmdLQQkx7Ws2N3W8/NyY1B5ET
xCHOaEqzpd4W7+Cb0yrwav6bgbwwPOHJcYbPWvc90KsQN/bFGj5rzMbhQfIaMoGr
bgqDgSvOY3m2C6d2FfgiHr6NmQbDHYQXX55EbsinHGIUJjODMqbLflp4GoIwYdne
ONzWabiZgrkdsYQpfInelxHj4G4p6wFHgHIoHyCsmvnIS1SAYxCaqYZyqZJf5VVc
ALHemA7SWE/TPlOuAtGB/fE8Pr99Z/SOw2I4qyk/a35xusmcZyuuYtvmkZd3VA32
CdfV2Ge9/jH/AJZLgFoyKB8CCm4kFZEm6ohvorURNK7yWZVNNPvrvaqjglLTHI4x
pT/7x/RqFLeoCOAvX9v+oBngHAtwNoHft7ZEmzJnLWaiBxBBliTia3A67xHpl1eL
dKv3ol32nvkzvIuRM7p4gsIfFLvEk6/aANavnvQ7L8iBJb+FMZKWBFoZ22H49xJe
hgQ4NvbwTr747ZNUTYv60lXNo9SHSrquBzvm+XsuOcUDeKX6hAtEl6SWXtX3PwtZ
ze3mVd6d/Ljv9iF1Vil57tHF+w6xcAarjx5U0SWNSjDSgxDdGfHBURQRGEUt7pDh
NeWpQAoOHMNIL9NWefJt1HUyza8UfbRlqorTrZuwNck0SgelG83DLiL1E7n//5qu
ly0w2RzBp20bSJA6VOSnRuTs1EnnxRMcnI6/Qtnh3iJ5LbVflMLi5zlU4rQl/+CW
tycNkSe6nX6gQzAMLjoU3Rsm83QtdlbjGLPPjMZqVRDoYLiOqjAkvYabdeG6fHF3
pTzVFMYsNxj1pYeBKiQL7NMtfKJow5V6Kf5r0XWjjwoJoV7Yyam3DyE/7hPEYyAv
7Ngy+ZO7XwpzerxHyWTSpA+Pj4DGjKrfat4+M67xpJD+L8Kos/4QEkiervYlDAjI
UseLxM+q2/NgkG2uTr++CJHyuMFBgNxcQ4PMkJpProXfzYubMV+gy7w8Vee3/Y/k
BfZQhSV9VwFuKmaECpSXU/uX+TnHL7NzIJRGO5V8zU2bxUTKRqOfxyl2orZsigQv
TiJA9sJMRXSUzts8v6KGyEVdN0KE1UshMeWR3VE1cTxDluIX4FOyfqfuYuK1hQBW
OAD9NDyHME4e8536CSJetC7KTOW5zYtwhX6m+US/fkJZWSr88ubu8Q9JCUuxcX3G
JNIicaSRNQ8iiL7vmRNFO5nor48S8sMj3GorUtHnGsah2YJdiSC8krRg+Twik5AB
bUBH+Hoo44NXUqUBAb59sfIrbmDwHNiWLhdIIfmXqSq8MA7zNPgpvJcHhiOdGV00
4M3q39qTwsebOmPxc8ffcA3RtWiOJKg9UiLrbLRzNhB71+cfiHKiiBxt5LvVbRjv
zwIys2YAKct+EXlrJe3CBaZHh+/8YSRj0/5P66XbfrW330auzpfGKIaIT0+WnnC/
BHJri8LNZ4ARurb7sHxcDMB6XEg6ys6KudMllicC7oD3ZKCc1Qlh/OVDP+Wxgxrw
siDDMnPEhQi2K531H0kXFfc8S0jdgLz7y41XbqLrXcssEb03EbaMhq0PjY73I33I
vBfchR0dHOmT39QqB0hvt8OKkbJVB+Y9ZVgvp+kUkMUBX+Dj24d78ZjLU5pdXJ0S
XzFCfOGWZCCWCBHCOnbecRSoApJV/oyU3u5GQKdpT3H7vGXipgZ+ik7MkiZbGUsy
ZhXmyWN9mFKegYxHjMffdoIDYSA8CPZmlQkt4svrjbygpIcS0evAthn9Vi+CDCEF
KJ9I8WT9oiBlh3aPKzqtNn07vj5l32knqNvSPP/DOurJaXyR1fY9MOYKfOflRSf0
h2DEj/Pv4v75HtIpfSe5ZnIQgrkEmVVhLhdPHsmPBBfviEG7EU5gOnXz212gQn6P
aAjSza42yFGy92/0tNTthjjPlU6FnLe7+N+k8yebbC3JZPfiMeVrYghfZD5mG0kQ
uFBAOusxb3hObv5jtkfDh7m6UdqQpFrkmZ/dP8CjNwFv7H9B+Lxwb43zQehATuz3
HYM8UTYS1z3bQaulf4vcaPr6sE8a/4xWksjgWyOiSP6sPbmVrcotwCWt2AGCx7yr
K3ZwnL/Hw4PvReYoB1XdurkzMpjgHzHkEpC1Ypir3DTGR1dbOeYvTRkFh3LgF1pa
x0Yl5WAvI21piu9Zgs7c07dABdBbWVqucp9YCVeO3u8VYpkpWMtHC4X5WRFTup/r
bQV6nlLh0LjfGY8rbSg28OiAtrODLlCOpz1kGA4nMbTGmaG7opaoHQfzBpu2wAjy
r7RSFMF9MPRIV+jbb/q3+8WFZlNcJ4u5WYRWOSJ5YRgtrCwrxkyAYd0mf6jeNptn
A2QiWa/F74KipDOQGWB0E8oIgXRWJXxXp8nOYi+UXy1moUeu0fGL6MZgGpFcQ4lw
XkNgW0a2ogUeSO58MvnVRJXW1eAlUyUb6O2KmDZjeBpTob4lopsV5lsO2UVgd+gJ
i/lpaKEbqiH4PemTA24VrMv27VuHJ8iedxbIyl49dxRqj/QWO6glx+LeTucPNoLu
BI3105SburS6ItwVnn0Y2zfyOaaFAmJENyJPMNEGhC2eu4c/h42op8zi461NsFNz
YMnzpb8H9dlfjDDD6LrleXxNA6OXq8bF2Y2QieoCHRnFqUvC7apw2SNxlE73W4B6
nTNEsg7hG0KC85wib9K0/p0IlEg3Dh964q6EbqIxqKr9uXDQRs7TC0rDR54QUlG4
KhJ5cqjDt+66bVeVX60I7RVUDkNFzVkQTjfKlYJUexwIh+gn3kHvpNbP1N0C1S4E
3x8misuRp0mUugeiEysC76tLYiuUtw+OOw6BpI0cpesyfDxiysu4WNS84d7OYssj
dbdStyl5OtH8+BrU/jATcrEK+FbYhd5w4Dpj+To7gIJ2bf+TVOeEPEuvswCY4TeW
965ZrT0eksXGO73rT70HLLRqUcnVCFs4WI5iKcsdo+GwNiG0DmSifbDKsQgwpJgP
0mDy7uPrNtiskFeJdMcDnMabfm6gCPJuG7l4j0EQvZIk6V3WCaQO7B81hl1RXIEZ
ny/R7QjW2GNJH1qA1nMZNKHwtkokf4tmpUyRCJS2mQhfkx4kn6GGmBArNBkjPHLT
4RlkXtEE7BMrwD2ND3m4re2C6UBAjRuFGOPR6MioOjO35EUa0ACBe4sZv7s9xFsp
PfdCDcW1krn9uig3rw6nhZe43yo1BFNBxP33vQRA1lv+Gs4NW3TzPRlXQtjr/3TU
hnD/vArP2pr4blo6UGGSwJQR4+D8EorBz8V++a5mNdXHqgnlOG98UFL62rEbTnFY
OK/pmLEyCQ3GyRovMvTFknnLTLp70YNtj37AAdVohObBcKwTV2CUT4h6PT+hH2mW
eTQ3ToG835hgM5Dqlq91/HUDgae25Yfcb4LiI8suE4v/W10VuNswtBxSvuOvUI8/
k2/xbYp2i/0TmJy75yxM024PHa+YBl+s2iz5iFXJH9AX5SqVp1n91R0Mh13VWu/V
ZRufNQJg6iQg0wIvrdWL8qfHIdqp9RJSybdvq8v6rZyzFXc0UUnesMW7CbIdkFTr
8IFEYiDYLwKLs0KCIR3nJn8xDiPlKcCCrk1oytMpFfGv6tZ447tRPPHKxVtfNpgm
vA8rFH4F6/xhcbcz4vQ896UrMRJNwZ0ZGXoiSyo+rf2+K/XxqDTLHs4hxS7rCX3e
N5Ca07+gZ9fyyzB3JiXprJXlLRAUtlgwpoMbyNf/fJZwiiQi990s4qw/xaMkOa0o
qF4tG0547rHs5IVGQg7mr/bKnalTsCikqPk9/7x6Ya8MoJnnAEN5h8fUJVM7iLIX
+7pyX9Pf7+i2XOQ+wGDFXnwTBygxGUAeCNb/WKr31vUqHJ9yAEIr4aTpos6h74Vq
DjSSNzxZq5dBu4koEyBHCJvpRGwET+KFRV1H1fTVWHmcz+WT3ZdxlmrrL4zVMSD6
dSIz13d/3uxANaP8RP2ZMowkhhfdf6+mYhetk/9ecwnB6QmRRtwV+krLrNq6Y+Rx
VVPpcDCHYjOtoSZOxFg1OJuixWgQwuxhCjGWl5FN9TpVGIA6GcRjfY6jPlpNUXYd
ISGN1wuJaI2NvEdoNRLeO/ShTdLa24iPJOektNi/F0982YexdSQngWt25ke0OMi+
mwurO0CcQ+/B+3Ds6GqsTQ5FncsWj3mGhvO7rELFB8mc3ucR5IDQNAKXkGkGea/n
iwz09NyTu8l+SLNoQHh7wT9fbliyQ1OZKT33ncKqRKv1LrRIAbdPPFp8go4UfGRr
gnor2X775HybZnw8xCTSb/jITJNwMqJ3QJouugQyymqTwh4lbr6cavzvCLhfizys
SlzVlNkGyeahGlI4E2easml6qent6F4WNY/8QZLQ7euvCZlnimS+BkGqRpBT/5le
fM7iYZCda2gNHAzd00xo6RXFiMfUpFIAAAFn28Z2M/mHb1JDmMCUVn2cFy5aWcuk
gQa90FLhsUNEjpZkJzb4fMKVoBDCfRKZ55nefKr7gZ7yapT7WeKMINYcT0waX6uQ
ULkno6fTNiW9Vp4pstSQHOajr2ATcm0gDSwe0fW3f78c0mIx8Tnto1nrXLS4L7LS
myDBFGsizvZDwD8wZamOEF4wpkW8K6TaCosvEnbg0eQ4yFxq6+KD2LOBnpUPUkFl
AyjudFV6NcfLze/68nqBjEj0WfUkmGpFm3rCRMUc5Zx/Eo5TOfHbjyJwgyxmGtNd
aLztm7BQlC97m6jM8mnP6lK+wW1Cb1bFs9KeqvwtTZFLpN6HYY5hVJ3bgyVEKg3w
I2g/PRSchQgZquDa5WZbtEx1mZSS49HGMLt5km36kiSyuqz5FtDLv7p3XJEOmWK+
SaXPJmOpcq0Xj0SwR7Grk/Vv69LnQziQ2j2HPnnUZZzP7zrCy2Zeey7U6GS6+o4W
UPmAusmyS4LL/54ATRL2fUUxeTvkSLLRUxBDpRO70WGmiE2IzGToOuSAMffjrNEx
ql8+tRAaPwteLWpBoxDetB2UrpitL1RcRlFYWliD3v7OCmbSt7Qoy4myDSTknYdv
d0SIT7KDqEkt9KYNd6V/8DTTO4iuaq5TEjz4zNdUlbJUOIq4iH7qEYqD3HKa9cjX
ZWxEbteW0E5056A/fTo2e34vreqNGRrS60xUzdS7AswQxmpZ/nt7IScJrR+HVLS7
bIJ7PYGXFBseZrYhbP6aws3wczLo1SuNTwkpqgzz1P1WaaHfHAMvI1oVlRTVZjwd
7sj4HOO4O7bGhhKoykfpFVqiXM260e1FhmpRdWUTqDniIuCk45ROdNmNH6Syrp6y
FYI1lX8TCqTecHLNk0LSr4ZHBHrNxcXK2PnMmsKkt4f06NVVGwE32/HZ639u/mRi
y1OJ5QNFWceyhYk5lPpvNw8i4ofpOzU2O2Zm+nnMD9zs3xg8leLaTnLFR0vlmi0g
JoI1toLT4yGb5axTnJBJfJ7kR8WTD9DQXWZxPOel4kck0Q0oJ/IOf62AIMUDsVLi
cFOEzVQaZgt3XL88JSFGzQ1hdtn0j4UWUypaLbMoGS04iIld3jxV3KGSWsp6HX13
gps19MQAMljpM2Tk9DhJkZqUkZI7g8o+ZRDKJQqAyRI61Ih6XYmzlQ9Co03tPP44
VoQ6FWBk8qvs3AEKItmOPZd+9U1qgxfRAyLV0uz/HJAqis2YTVgZ7YeYdRbbdwz3
/d7Uc9MsoHOHZpRAhZLbpz7RJSp46IzrfHVvJjsx9vuJaVM/XVwB8WLuZFT2UyX7
3cUimztYwzzeDoHxM5/zMhA3ura2vS3urnWFw+fwEUegvqTezhcmxerrz55ZRL+T
DqMWzLTY3G0vNF5E9+XdYXD71H+m5B2cOKrgBKCIZqq//2KPw6z87bMFgyZbJ02K
4ZUUSie9PbaqES3DCK9WGiwTa5o44SpJg7em45JFBslT/wgUfzGKZVpqOi9wgfst
SvV1irm2wK/YwsWUF0sdhNIaQ/wIMqHz9v8vHLRlczlUKKth73SGQxqxmjk6RFiP
vP2pi8LbxVY3vTISUSG21ub/oPt8Seb+PlnN5tiCXrlkHuZb8juhwA2KxX9LUE0K
Ffy+QRvME0sUQmNo01KV9kfS6NiYtKG2Ib+NFmK9hYYfTzwAg2GOvneVwwfka1XM
GUsCxlcABgebL5jH0ucQggCPVtCq7wfipsvhMh1Lho4Z79OAgrbCwa9tFzdkJSJJ
zQqu04sGzria/uSTVgc58FnVm9+hspCQ9ziQOWa/8A1YvvrvXok8FrrMP7pCNXPH
jzgrhRo05k2bCyEej1mVCzMLR23SjCwJtp+N2gkqVsRp4KGPJIY9ZljrtrGpLwjB
XrIJK3jbElJUVXY8iRgI49quPdk8defu20coecCvFPR/uudwDdO9Erh0ouGQEs4+
q1eHujg3hqq58smVcDQscWHO6K9dWex8jgPnnaJj3lAvr4DgY3YrG95dWWPkR9W+
8hwLouwJQDMKvo+EFAqQKeVrsUFfmQhbYsG5GocTcUFZNmM6tDyqWJ1BupC7jyxR
xux239/Kj6Bv+CiR2HKOHmZmqQNCHSTNL5yHLAkAEFLzF5QHW/TPn0zKkgz8laEb
5DhrZ+9/h8s3ehiKvFjGBQn22votgNKlZbXSoUyD5RfmDcrCQxK2kqhJ6y0xcz5u
RH2MzYI6rsHzxycBfLNhRlxj6SycSNrXjAyX6Lr+Gha78veHoon5YLpwEhSROAcS
WFa5Ke6RF50hB7EyKfOzs2SqAInGp3Zy7CpuTis2fQ2jNCQUOvN8/q+jCD608zP/
hYYVIsZdQNz84VMFxXVO+5WjSN+/hN91EJMa6D6A1m2wQglBPSuelemqVgySuhKl
NBtgyyMsX3EDmDt9fMTTolcGIG4NdhLRxk5WeROZrUYn3s3gqFkCrFR9HbRoC3jj
qhFbV3C2OlZy+2aO7u8OVBAk9rQPiZz+sXoTMU7oMSLhNH8o7spG54fnIVDkHRVC
O1OjEZpI8WNeoJ5agIlQXA1SUT5u6r8pPsyZNIhEqviksGERKl1sVOJFDWxAYblJ
8mAUZCZpWHMSL29SVWD1uxBa8mKxNGobCouxuk+ooiDj7WazmzRzxr4l/TuJ++jH
nUq3hTs2QD6euvl2Vv/fY3sOUuCLnhaDx38R2k9L6hr8XfjRbsvJiFjOPslxfFYL
P3137WmD/ynVpn4hi7BVQnSkU4vVv2nNEav88hfZdRzCu3KxaQxpoXxK3lBaP0ma
j1m1XoZA/MlVry3K/phN/5qzUjGH8RXbSoZgewCTUXCnwBiy2KN/Sx51DMqhJMvS
hvh7cgZVQbnEDC8/QMtN2nAt15UBZ9VxLR2Xa6UNUJi9MQTDY4NcmVPhus8yNmue
XAg5XlOy+9hUZWJSd8cSnVU+++1PiMHLGv5nfcacB0IJyuwaGXTrKa6U7RzIPQ6a
jZ5M1K6YTlLvimxpSmedJgjdgER6oSN3HG5Q1H/u6cqrsDlprUJc6upIZxPNO72v
buBEoNGax1RmjTsK0cSfFjgbJqSr1pOZD96llSi6tNgh5KZLQN6s2dHU1R3lTz6Y
FFZ0XGEtK0eoqfokWpJPFjx7WmIm8JilzCq6nF7fbR4pE02gYQwFOHcyQcUnX2yc
IdkjvrREjIFK2XLdmFY7xTyt8urCa+ICW2jXZdqLw43p8+JI88PWeBSrfg4MHmlv
wO+PdI0v+jWu1HaRbKAV4pPRoKHtsDwBeMSu8CAp+kf+Ae836siaVW0IyPclP41y
2JICNts8vm9S104GRVfoPV+gXELqq91dmDcc919yT38YPT5F06CQuInxQWVit2xh
xU8+264meTozLvILFhUCljXvcl2HhY2GWkUCk+6LChw6ASjQvOKS5VreJGCo6ekb
LJeNZmivtYJZeMNFga6Ea2tozqjETtb4y53tUS9KsITyZoQ0jIFqUtaK7lbPuVCx
C1keY9q0vCDC16+B+WQFo9kMOOGibqYPd0cnY5U7MjNHC99MNayJib8gNrZU9BuI
kWKyXQFNDnsXReqjEh0JXytGsKV9jVmbYkmx/BSjsWWSOdl3lSDIMfMOg2alYRad
4y7W8gsq1umTb62gEM6rmuL1Se9O0OEfOQQmWq8oMyS49YZlOExLstuu/HLq6cwH
H3zBw0FF4J/tIuXVQcBQ2KX2DSgzhe/3epfUpJVtOIKN84yJjr9M5UHXvaiIQzTg
HWEiEZxqt+CVRZ6fYrRX32+3QdG+RbmDCu2uA9UisID8cGZevL01kNZRCVWtWSMZ
ItQJouenKTdB5cAMR2auakbibea0I1VqXuE18vPeEtjY+ibfwvxfrwq3ryvzQrxP
IdAOggxG9i5LvgYo/bSkcJ40GH2ncwlIOoz6I4W47BmQ0ATzZdZ/3tRSGmE9yRtc
AyeIgGUOYdb6XKu8D9fsCLykk9ARn/V3iWQrs1vouE0elbip5ar/nefpy5a27ZMq
dI6LNCt+i6snQXPGoWokNyZ979vVROXOGS9sQfdG3Jo6fxnsqk5lIVyrt+IESK17
1Mm2GV+CDm2xIMQBr+c8cVMC57gg1q+yIuEpbD9B75YFpNvIz1kF3/SRP/K8nDM9
FTK+oONgcRfJssiluz8m/PT5c5fnHklGWxAD2+MT+pdXYD5m4JmN8FaAMp0bwXLd
eKkNQfyZra742Hn24NzJN3GtD8P3palD5N0RHg4aHtAXjc63pzp3rIhly1zDwDqq
EygOTpeu4j0X4MNxgAueYFmvkNSk+gblPe0d2p8SioBR6Sh/HpM02V27gOk2+5KI
3WzKfEaymTSEjQy0vw8VIELLmP6lVhCX4pCaqb7BqSDj+/85l2Hjy8KKGNr6ZJAl
lzrqLYMy1i46UDHOBhCs1m2AV7uHoaCq9HAvNr8RpRSEYBHdL681+sTaThuM57gJ
2yFYAPx+BOFKKbnwywDw1n+OoIw+Uk83ih6Uz7ufqDvyMuyvwdTWx2AFr3lj0Q6g
P19Zm6vSddZqo0aW4aqap5BKaR6jIZaextkONdlbObPu8Gh4pDNUtsczdajXWPnP
6plLsGCp3SUm/qKAJmp1gp1M0vMKMoQ8czSGkmdrnZisD92jdWd2lCWTbRUpDQ/0
eTDTnFYuwXUMCGD8GRwejatltAjl7SKb5mGCPyD8uHJ2JnJhNK0JSrV4KYofIn1J
cWUEvsjpVU2v2Msoyjhj04R+5GQGKLrD1RtV4cBIvxocOS5g5NTvQODEfVy2EXuS
3lvw4Y6h7FVpRsnJbhpxl1YWguZ4HWuVrKsxa9ZUTWvuArfYGeHNBM0SHbUOraT3
LxUkJ9BwMFneKBjqBcdhRomYielWe0kW3DaDAYe9nbfFs8RpL7vfG4EWtsKzG7Pe
PPU0MoXQ8SZBW0tWI+UrY6nGCaDCGcjiEstoqKrpAYpYG4rtnqIRGxk7VacUNwHy
g4Gk3mqh4dpefbg7HXUwHPeaASLFz0ulLPAeXIC+2reGCfASacm4Z6zajUgqTT3s
HOnXrTTVPeaDhZ/qFhzZDC8bTnxE2Zh7sThR+QwRoNObvFCNdVUONca6+VjT1oh6
kAYOeXQ+FGi2poV1fpkyRvFpuNwAecJCkxLRJNZ1GUGS7TxZsaBJiA2QbKklCjZl
Jkg3Xj8rTTFbMmHwjBglZXfTLps3jwyOyo11pBnmt1+eKU7gbTvA7g2Wl1RjzAv1
9vig85qZy3zPoZ3iF+8+5uppto11IifRHgJg3kD10HWCrEzCWNgLWg0tGKk2s1MO
fM7I9Xw0aw1tBafJRtEGL/EWLKaK/WjmdBBWdiKf1tOeOuaIMrjTVHPU8iQtQX8S
/xKroXOpcu2X1FRq+kf0Rk/3Mzfug3/3SEB+ogUQ9JJKlR1fG/GrQHbKCqJFeLC9
EBvMG92QYu6OewqX/fOnUsNw/PPAZqtoXBoUZgiL8CY+btuw/JOJ6NGT6C8AGVHS
4QsQPju2rPLSPp/gWg8Wge0DNAiwz8Z2MbCRP24/YUwOLWZRpOpRnszcCj+Ck7Eq
po2pgkuL9+amwOxZOB/xs2/8fdG0FfAvWBAz0FiXf5sJkbVZy6h9zuXfkTqLxh9Y
ZbuAcTGLL+Yw+CVgUioM6SuuCh+VcIM6KrwsGgpYQsn3z9FMBew0LaWIkCtxF7kh
fPkYm3IeM8hnFxeMOqW4UFCwqyWJ0iczBB/7Lp04NzB5bfaGdxalkqFRdssvc5fV
a9Doqv5YDz96SnMpijATil9dCZ/V68OvClO3SSPlxb4HnsEDOxuJ9N5CGA5/Kxdy
0kUKni6tOPqgAA1OIzvxKJws4JQRFvcLK7Z22GN3i90heCVylaTLk7KCRhUWPu/I
7+lnCHmQxuO5LcuGu1TVquyTjtQ+2KDqT+DOGT8QqMNQ9gapQ3KpT/SMdu0L/jYa
DdyRbqoibwqdWgoKJHprMVHCdX3m26yEoB/lvllCGEddlMg/Hh2hXqZED6UP07kq
n+0Tr5+R1/GsKl/mPYqJcr4dQxFY6XjaQ7uaMVgrOnLS8hKfePeCUm9CH4QT6MYf
vsc6ps/bNr9QGt+DSWm4klK5SrQTeYmvapzJ790sSHP0MD+RnQHXFk6vL7Tz3310
5+48Mh3vsXt8rM0Oo4Vs/l8LX+O8akyfb2+4iqx8/dPTMfp2J0bG5XgCbu7jPF8y
UWXwtqiLwqv/GB0C2JuOC099NXHW3spdHxwjoF07dl6ay5JbcpxOAS+5FtFuP+Yf
BdKZZW0rp0cincqsvHvXvuh2HPYA9oj0YEEEszoOR68/HrY1LwXBEScTt0Kl9PuM
GrXI36SbAT8ioPmF4Vt4WTeFRKi3oMtaU5lzfdLGrj+tT19nqqRL8eI4mQ+7nuER
vtoJBO1aNKXGyXatK578kb8XYexdkUfO89PT6OSF08g69omkQSwJSw7ft1AmuPgW
7iO4wiNlLsJbeH9obA4YdGdIJdpJbHk1hLOBaV6q9k6j1SE7zyIJJnFTu+H9Ewkl
HlisHaO1R5IWLAFqNj4Q4bVnE8Qqc/EsBBhaSuTN4IHbfMKG4Id/xNj/nL4NxvBw
hZSlEJk+bwMmRdXrsioMtlEZwU3dlje/MBUmM7BBzn2tdOc4LxGRGLWtRMZxx+5l
WXLPc2+jn0qyk51lRr6phBROqUFAiUKEMsbIQsll+Xq5mOjs0Y33bfa/Bs7p6OCn
ZPCtKDajVJnlUDmNqLwRU4yU0zqoquHy58fyzQT/pRusBYaGp5JLEm+6HDkGQNB9
Efye5NGCCfttslvhKyjVTKskUd1OrnBiDSppkHOE8SSA66EFsyF7tJZH1m46ngb0
fVUYKouznVhEgY6/IU1HGHgQRe205Db+tfRcPciAmUL0LPv89kUBHEKKq7qmXjZO
VQ1UCTV6+khnB+NgysFi0QLRC9Ye2/zHVqIHpqAlsK6Kiq/M8Cs6WlRQL/hzLgYk
qkuGoCKLz/KhCY26hRLaMk+k9UzuyXB+PMgJXPi1KcBEEJyVBgj2a9pk+47PbvP0
biB/ZXYFaWnpeZMlPhlA+IbZ66rTSicCzlQ+Ss6FMCn19Afqj+VIeicUyt5I/9W+
i3vji908+VXXjn3px38768iEhwPia8k3W6nTSG6FdUh0VC9jrVCQYFq1f+Qz3llp
4brSArp049WGQWHCfKKKppkgJJIyqlpEQSoZHtqnh3d/b+0sBjTXZSy/Nc0OYWfn
4zE9Wv1oyEzK9clliI4FeQwaHgyX0nxioDT67EGLwQCTNzYhyLJh0w8jAagkP+1z
/fGrLaVJP0odWrTZl62iQOD6o2176QlRUgHCQICr4u98v8VtquCAEyXyWFrN9dWs
SyymNGcTUYPydHOXggh3eB6ZSb/64X9fx1QkWk1Knp6HG5mfCAmA2csZbGgcgOik
ihHpOZ1zQSEpG+KTFCjLE1hOvtb3gopjF/fTuwaFEfibIQgPk7JkRZkRTHoina6m
oOnZNVZHV0LoP784hVv3VwAUI7FpTxKEgaG65/FHvgzZ063MjDVxd+rLqyF6eG7Q
l+s9mAI6u8AEAkI3TNQDZk2Hjj5WW9C0e+eh0ltJs/3fsXZjfTU3LGvHeFXyzw0c
OadoKT78yKA9St//c1ixjhfl5Bbzp7kMwRsm9axffNCWrTeZch2hcdT6axkL2dGm
6GawGHX/yGGNSLpZAKxzIpWQjIzbkotBHCBgFM1fkcczu6zbtMSUA6mT0LM0jgAV
OMUS4ls1QgMlmku2LFM6h+65S0jb9FFVTD5GCVPBwKzQ2TJot2ZUIDdRFeTZclv9
WJsZQNwgz0qyHooVtxNl23yTGDza2jdFtLjcyQZ0XwHunznS6FwsvhabUkdS+ttP
5Bbn1YJFatcd9CPg1lQ+tWSxQJPLLz8uvN5jO5/BRr7juNBLm43dfocS/QPqJWEr
i2qbRGBDQSufB6yfkI5sfZ0P5RwsRJAHTD4ZlQuQNqVy1YJ9Zlv94sU9bT+MTHiZ
dA3xtzQDJ0l1yaO9+tEwtWbe/yP07jnCgjUDaM2KlaZgnib/NQS4kxstwhUW0TfE
eAao6654MATmvQQzdE151Kayxpyl0/z5SyblAtYxzzZnVDpUFmEGzycjaurn4Dvm
vhpEw5E71ug3HEy5Km+9R3RaufLGS3ziUJ30SnvHFheuJM5gsmeD/fQxtBXllsRE
NBqiNTS1TGOh0pt3Mo8gWi2uL6WNNVoA+EXeIulo2FLbX0a2gfGDwbiP8Yu2SFyS
3UAcTON3DJ84pHcUvD3sL54+gSGPH2rQAYBDSbevH0ow/S8aK3gyNoBlwzSWRBjr
jhPsq0rG7L68k8cgyYOifXHVz/X8QmJiuJzhbxBC4artUDg/7jLcb1bIN/MQ2Mpz
Ksat+wUriZgnvF9cZ67nulg1lfC+eBj/HHjKM/rEEOP6ffJqIiLeZDALGJrSulWu
iRIQLRs/i91Y8AZPcw3HFS1fPtzGKAc28J00BZ3ahK5MzffgWn5S85h4ZdJqdMa9
knlQlLfRco0SRJ6BzEKoBY/eNwdaIEpVVogIo53orxUrDfe96C0BtfeQOijEP6I3
S6S3mlvzMAgSDvEKCZS4yhnp/79uushLzmGLkhyReLyqMy7P8TJhvFGkHcYP8qYa
lKkjQ7nRibiZbdwh2Zx2FtdFiOPT6BTWMoJNbxrTcH3I18SgAfJv0+b2vecIFNH2
/fh29lGXJLB3JxhBToh5o7f0yCszrFTYWs8FUgHB4+l4vRdy/hxzlMu9mjDDpctb
sVFunEYTCmPX5y39FatOT/DMq3bzsDIjpbVm2OD1TYULi/VLB9fUF1hN+ehPt5Us
XCWcE+a2IoemKyTmac7VH8OtqCKxveygfX0x/NjGaqTRDDezFb73UZ09L9CL26en
g6tQNkMRvDKCK/Fa13oitjibRcwiT6tXWtfX1na/jLpvqVomD4UbzsyjLUGgHpxZ
GSJR4+chBOXCFBXseDCgu27vVv3wKkBdNW7aCUbgxdl2tnXTgb+c3RQUcLeVAzyk
0wmpjMylX7ATk8AQHWKFs8lMIFYpmMe0YMhj9aqbksyb4hQi2H/LkTFxe7HWmzOr
zfyBO3NJIM5k/wdDup+vdSkXm7c4JrWUQX0w4Kp5E9kTHbeh3T8KNWbi8b8zqVNq
MiTNn7mRloRm34K4MIAzHbTpl02CpDsXpcGuDiW900M82mxgs+Fixkoi3nl8PeyV
wo5xWPgHJMC/BYpm6gopmnVPvNFtqLdvHGOhC4ELcJWp6csIopmWu6alJ0QviNwk
FSj+yQJLoyKpIJxv8XM2TvmHDk3NNW6uK5/2axE+RalyGedZUTBxGTi+isuz79B8
eGqquEgkQKxfk1voDJxki8omRV2QnxIJrdtZn1JF3B2l8KldyFDZ9GW8rQc2bSIo
JMCLqcivCw6WjaFIlxBaR8Z2s8ejuXFAIzLrUY7CFZZyNirDTU3LmKoXpIKFNLyI
Vs2/gaDHsOq1MOmUeXmAbgTDdmEyjn8lQPbhQCsa37SU5EUo7mrX9LTQGuVVvNV0
qqm46p2BbhEmEdIVb+zppUhpkKFBU31zKFSrjhJ4CBTIJq2m+k7roQ/zxBnSZ6tM
0R3SYNp+txyL745YXcKNOXE3fJA67u8CHIKW3DcWpQeWDFL46B9zig6itHjzccXP
XXAGAsIpo3ds2+0twqCJjucs4VJl7UHkWKaQkqrY2gofO17gZWOXWhzvmUGXjHnG
DCfma62Bov0Lc2TYYtkWaszjh33ChcLF+vDlg7fXW/9yRsSO8kvgDK7Ks6odk03X
MeQJqTA8boE+3km9fse5U4RPtjtyY6OCYmoUtWnqBjWnKtQVdOj3BU92cBAMUtwE
ceu5pc8UFmp8RkOzYeTJhBiqTp5H9EsnsetKWPOdJ9eKFkBkF7ARefltd/dO6SyK
HjE2+oKdY0KTRuJMQqi48v8Ho7g8wvC2U0ZmfLEMRZzTe9Qz08uC60elXoeMSRwX
dXCVVzJOmMRl29A9Lf+/PDfGHm2Zxo650K31LXrFYFb9LKIbrreCZLqOdFUFZMl4
HEfrCObGmmcCAIFFupFDlZ8MHV6oCh4OJjqEdl4fgx/42bFa3oSIrODy6ZbsXpqJ
rqbz/bcOIxC4yHDgUR7HqJB7BoE0JQENe0xUITvEFM0x18ezQPPzpoyZ6RUiXGm0
1Hczr7c0ei2msU+LR/oFdyU0gLH4mxhbqC04ah5rs6pB4eQQ3030R4/olzJBSBsQ
c+/rOwScwhULA9ao1cQOb7aljhS3HGvd0ewPUfPiIehz+UOqQlkXw56k3gCeKrWe
6blBFHttaMQRh9f7joYESrh+m8/F0ZaoELLnhU2Dh9XGXY7GWvuzrrUA1g8tzoen
uqZODcRkAaT7r22fQOJk1pF0aVokeD6EzdI6d8vt444l2MGRcH3GfjoaLwiGjWPj
mG3nUr/btFrQmIhQiW9z1O3BKUDq0NnIPoHIDJkoDW/WdZZPUKYAEGjUCSvoMzRM
iplp6Ho9BRufMLjyoOhnwUJ2rHPKVqABUqgf0Bl2Ur13QurdhwFXR6mP275qWC4j
nRmrs7YRI/DVSh9CyJh8Nn3K/w+YR8784HlAHF4D3It9sRtb30lbheu/EkYVrLbS
t3ofb3tMRYNeRZbUoDf+4OpW6woBprxkk8qWmlmXxr1c6MV5IzMCPbihFcBurhQ1
Qr9bko9t6MwjDcDtKsyJGNMzv8HcjNs5Kg0O8E+K6TmJe/5ENxvfvJkCmlUWoImP
vvdTt0GSUtomikZbcIPhEF7FbuW8g6u7BZNMVGuMxo9/HNQgVsFlxDrW71jY/mfV
/DLZqRYpsKmFqpUP4/GoFpnjmyat4+pnngFTrLVIn1iA3UiwFWcYpq9W2VwSW2Gn
lrFu2za5TEdxA3ycZSEH//WIrZHbc5JXfXbJlUfAgh8sAqzAMeYn42caqqBvOe/7
QH0ME2TWrt1dMOnjbPXlLz3/YyUk4k22BHQR7Ps3Gn1WD1d49ViLsxIIQ/N7AzA9
YdG3AP1ke31lKEU2FsYj8JRYo3MjXbvyWCPxNFMJR1Mf5it5/C61YOmRb6rttLcf
fdTO6EPC3XTQNNoFsRaxWCC2fPb0EF0lUXz9SIE3r3KK7CkEStsj6u/kjRzRqzl+
WskWmMRXAyQ32Of6Fd8hmXNgsohDBG7exfv8zHCchFSWjrcpErwO2yUuFYrSI0KA
xDxvc5rgQ1gTrflmlT/azqO+4oDuBhXUgeThoTop/L/xvnCtiA/5fxvZnTn28XwA
V0GPykl7XvyJPjOhO4ICP07ih8COZnOhdR94vjVWKYbcpTP3LDatlWPV17TWjFhv
qegHrlzoZVfs46s0UAyH9VgtLAEN78LGPt5YJP069cSUX3B0MqvdwDY+tjBC/7lP
49421lX4jIGUoLs09zF+WtSUsZz0Kn5GbI6F9vrMkTdHdX0PPxVgcQWcO+p6wP+8
iQTkDBx+lBFnxjtoA7vjPIAWN+36RznTyBxY8rrhIigu5kAmQqI79jJY0MrmQXYO
hXZUS5DHVvaS0SH8ooePjtRNuawBnMFSLvUV1y6tJF5zurJP8RqA4VuVCkU5RHv5
zeHuCYXnLLRpD11ko+D2BmLvMLfscORx/+cor8kwretLZ6duGnruLoTtWd56MYkR
TyCcCuinyrZ5vFeKarsrmeHVDeCCgPviHLWAuA8tNlOMe0HZtKRQogmn9rSLU1YJ
zwcLzcov34X/evSRRn0HoBIqUm2RwZ2PVmy7C8zoC1feR44EJXTPSaDnPjptfReQ
Ujips9eo5NulJUg5Ph3CUe67i8omeWOQII1oHUY1dYS1impwSFr/pnFvyYmf+fPD
qjfbK23oOhKCbK1vI61tGCx1KrAlb0Xwqt06kdyc273artFWZht3od5gq0qaIvbE
ygf0evPVaJ56J+p4xZwgaKJQzNEHDqlUV3RuxejCBvdMuv0+ZOqiTSoXdrs/yXua
UFHfBZVUZxUmFy3rlPYsz1FXAlw6atqxmHJwxlbLYZieXHBwtWTSR3VK7qBk2BnY
9j57kadH45kQKJcEODzX9HmF43QFMUlE9DuyV5LVgLRgpYnNxNydbwwR5+jO5hAx
9OvfQ6axjDJN3/FTIY/hdAEbXEWyTZU2CYwj+k70jCse1jDAq86SIXnGFP2Q1ZHo
UqXA7uX45xF9XZAH83glz1tV6VuXNy8J6ZdkwwJ5ruupkcO/JcLKkStXjt3e5Qeg
FBclQwI7+my60s4jF3aIkEpMkdBTXY5jFbz8Az8Frhd2CTwhDnhPeXzYcLbVgZwG
gfSCEXA25oE0lJICV81NW6hTvmzheEDIfwECcYEI39r6FrJ+x1+szuHa+EErVJ8h
QbI1scN8S/t525p5VZvQSeWG/8gt/st15/PTKvxxTax9jeADwvFAseaBbe2fUnpC
7H5vCO0LMLtZKbEYkRS4ljZ7/ENE/yQo4fYgyf/Nyem0dud30EipqelHHpmHdozs
hGRrN8DX2DJTr4GXMTdgzWSPcvz/Pp1Ia+VgH76lpg6gPzXi8pJzUprXz37p+JJk
yzDyhDcekMtIYYDL91y5igmu0wk/vszZpReuTiGntIeGvZOCoISqhX+/zlE9Xsln
SuJkepLDUoNklDixh2eq1NildGv9eA15iQisnIb+8GIK15vofDtgHDTJFVjfm84a
Fp31F0rVRKY6fRZ32yX5XETdBWGPEiytuoXlgkgrb9nvfEjh8X/fhak1RQANon6r
z5EVYaKumb42PuNnFTfio/incqqVgQXecCiSLSBA2cwI/7Cy64iqzDhyMpf0TH0H
LUHNMO3EHg2blWYBjW8IQazWlQNDwb5wXncRcuDgPQuB0rHQiIlVNOmnszFXfJXY
dCn+Jd+L4a/wdFnJo7JSeMKivknRTnRhRIHbi65UYs469P1278WZxxf9We8hE8lL
YRDrriMNLSJdTjw67IoLOLNzwvZ+g30onowBorI4Z2uF8mwFcqAXIgZ+2ePOIXod
Re8WceD3C42Kgi8TKlyW2Qez1NsxEj14UGhb8DCdb2UpYOzP9vDX/WaGOLykAWGc
cnEtTXyC+kxAHyZ5FyIz7KYZP9K0OFF7fR+gLWRq+hVYk2WyqEUKA19900uZR/0Z
GNgpwbkFEX4eru8n5BjiD7btwNhCHfKL9tyWDUnCYlKUfljijNHwnKdNJbnqaFl0
ZKmLCkBn6vP8aa//Eyzl+B7DDN7EzVi2zZnKcTRcLmlDNo9BVWL6RIKGmGWnI1Kt
PZxHOQI8Yj7Gu6/qkHoBV7PoC2lrA79t6JjQ994n5Wu2YRRgtS3MeAz7chUbXM15
s4bBtxYcITZndO6iQGrrVeOmZyg5Ceg+TTz+/nkw8lv2hgFgJb2tJ+9twuqFKQ13
QzSWWP9ajP/IFiZDTfG8XRjIPHitRG6pi8RW8tWdB/OdPWHnb0Pv8KbSoS4SkzXt
XLrcaq2dunrQhbtDoY4FeqL9LKCJ9qiS6oKSuOkXeE7Ovy/YJtMp/8B7S79zQeCK
+6M65OYs1++b9lMW4UDOE3DxTKMbMzv5RB5k7GK6La05eHJKb1uRuooowr+upY0X
H78dIl78JmAp2akzNGXJ/v70HI3IFCdl+0V6DtVFeONcLtbITpztLdETj74x62Ln
by95CHrHU7WAQMND0uf+3I49+AuSXlbCIlqQATgQALQynjl6VD0N6AudUQOZs3Kc
EnoAoBVRXoai6qgyA77px1tZHmej+9d8Ds7BDuoZkzCLhDjBJ1/MVP4QuI22/L/V
4yTnxr9io2snLORb0R6S51kHCz468ZwiCgm001+sqze/rtCxXt//7gOANqmcF22L
V1B+cA6laJcUjgLF9R0j77ZUSrTPUqIL8MaxZ5VLu3LDXIrXjI/AEmjgrSwzbSlW
GTAv0L2t1C1L845D6CX9bXj0XEGCsfR49Xrre/52hru6anpLk3AG3yA/6d3Ry3iZ
AFovXMzr451KQAuASMeJes0DdDKBLkv7v/Y235Sk9QZBVkekve/BB8SA0fWKUQTv
z0CBpZI6JHJGmDToksWzlGl4PCEcr1D9MXpM7UHCLA8cc8azE/XPexwo5Vb3JKiD
RYbjT8r+OFrBA54lfp4BOt/mKFu+QSU4+sJv0W9ankTmga9moUCENEwIhptRPZIL
oUi83kAnmRIDO41WfeoFeym8DGlvd8fqNXGZtLO1fxbaNOKlfr7V/3OUzQXhs4UQ
qF6KWKYKWkGhGWdKxStxbXAtqdgq1NCYMc+YyOTJAZ28Qyyd7csIPw3L/x2LpWoW
/r+tDyOHGxunrf1nB4OBTgXP0yluR1DmUhwSjV2HGzXC0aml56xZLzYRUNAVQXEF
7N5rE8xenTtuodKlg9e1GJZYAEkqWAjYm0twAax5aDC5pdy5YUkaruLgLXrsaPV0
kd2lux899bpu4HVaZ3L0UVUZL0Wn3BMy7vCWMClgu47hiODgsg+V3F+B2vOoxj5L
TjQLkeMDxitFfjuKfC30M6hSFKZFI0Idu3l67kbBa7o/BzTfrElUhmbQrKxfK9rm
nN7SGx6STB12mD+bt95cRtWzIzixWomOg7zFyu7HXQYDKZkF4PHMTNyKEXwQ3N//
FXc1giRuZuPKHgTjYu57ZCJbm5Z8381l+vEV4BzZO6O7AZTadFTFDGh2s8EeiBI0
dW6138DwZHVcBGdqwrpZ8PpnDtX7LtRxNXX0mZX1ImLXZ52bbfCKjk2ULydf0z+l
zgsM7P4U5fElN5yjbKfrLd93m46XHSvHRg9qYTbXAIIPXzJ3ULepJy1eg6PFD+/d
mEP4wj0xgVW20dS1fxRZ+aVSVMjrmJAj4vE+PKz0smzx5DiXDBoltzKACgTWx5tp
7OTRK4a6T6bha5tduuL4jWatNlD1klVhCp9XXDt9rALINhdupHGMXseiynSvlSyD
A2e1gUXRuP8KzCgrvbmktlek4KermgJsUF40Dm2E5cLdKDKAhRv5tlqQPx9SdbjG
riyS7UEQ6QdyAvVg+dvymjsfWbSjyxPg2omQOBlcG1tAytoCM2F9Kyri8cQC4E97
3scXuDqm2dQVzyIQ4fpSc+aUuiWjokZs8xDfq4w4j4NvJ5CSOh3dSw6Ef6WqAWCG
ormuy6NY4qyjkhdc3soIU+weYddVUimbT75bEHNd+n3iKFiZiap7AeLLs/Oq6mGS
DcFNkbVOKLAJPM8I69qzgX04F5qsst5ON0g79cru/98BINIj471OwyRj58QiyBXS
hwPPIF2AhWDe30I6X/NdDnA8X3cmb4O+Cx6zR46sYXNZDEMvdae8jg75xO9IPPgO
Xyh5WKmlBhellzJC4gF/cnHhAbazv8ug7hdLmDTZkV5XRPGTV3eTe+1gspHJgFdE
oW5pugC9Nduq6emdENA6SRmlK6Mgb2V5IpKEV9jstES0qwSZ03F7KLnLSJgKGRhX
k5uRt9TyhKbsUaZB2ckBDNA3ryoRGeYHMRWZGxppLyBPg2hBcnN21c/OZ1uAzX3L
aURH57qqOtc8UG17zrXJ4gfIG2wJo8wbFhl9GVE3n4ZtM0p6VMAKF8GqiAHTY2y2
WGoGSNBP0/rTf/RqUs26fNZAJoGmGN+1V+rrrayOHMief/mKvptv/Newby+9otNP
s75pXFPjA0I+tgS7SajdYaQt5laK6GFXZ6pvQ2CFsBVdcNRVgwD01N97xfey/zRH
6YmrivQXlrvYaMvaz6ECoe65m6AM/LY+CIWP6Xn/U0bbklPtdil5VSjwthgIkoz7
L4sbJCNaqxrhE5aCsUdiYx69jPYq51HoFgwYtPU1yLz8haRu5tAYPnA6vsjO9RwI
h0tWb+yLUo0vx3ZD934lUEceImxjPR4jAx3qL9ENvG6/iGGmJB/pLHJi6J+aebFf
9H9TTJTzLjwnx0ChapUySaBDFyml3/jmAmnymZALnwMTKeXAZMROD8UZ6p4nQ8Hf
brBk9tzqkEPkPbH+wenZVs5oIoS5j7TiHaKMepFpODjWETWsZy2iYsyeDDZgn4TS
C/seIpzEljNUwT8hImNA6LMDqDd1TMEh0ax1RL18EeuR7OkIBN+cYceBMTvk8IMO
frfqJiaP1lT2iGau1w787YxfBuVHdLbT+6Ams3VqZQ4Q5KyTIWtMRGirr00XbFqb
Lg3TIIWOaP/Hf1xywtOEyYChP+YEtf9mcw4kTzPVZAKVSDCTNNwbskQ/AV2m0GS/
ozxetOblef3WhIyS3e675hD86fXbLdq7RANcQv0X1Ws9h57MQflXxsOOzEXzPS9/
rcToq34uWU/r001XBGKNBxdhRNhY1WqiErWcu+6GhLetP9xGYMO84CGco0niY9nr
2XMUmNPbYIjaFhuAwTRRm9JZIGunlfKcSy31+kMxLx4cWk6PqD+dquTuRPTvqpGu
MbooeiQgBMN0SWyAPRwM0KeU9uwBk0VPk7/5aWFuwkrisS41dT80QzzfOO/Kux+1
4wn+v58W0H+CLJ4jWFGVcQ3XODAJy7ipdK7VpTZBq9DJZCCXPv4dAU9efNXclJZE
3oy9Ze7MCxiM4W+/8xOafQqdM1JTyqDWoGYbJEw115uWXA5iBjkFtrp3UDg81MYA
3CKyujYexj1hEnRCdjmFVfi7Rdgt+/wUN3IRTJq/TOcYHoydcbqwsnj1uo3kV/WY
C0y7kMgHtMSVj4j8bJVkujnkXJVXoZ1mMKVbv0eRT1eKXm2wuEYH9HEUWElY0sks
dqZRYcnZtEho1q6ebvK+0+XQicJI8n9WhfQjfVj9a1s1xhfBY5rUXRaHok1Q2tcN
6QBdOfYrZRRCvUGibGrHxSebxm1VoKphbmbmrf3lPn7qeD3qAzdqc7HEgRefJrhx
ueXMNxh2eVuwsEwxDBAGL7KfV9N28wcj1zlrc4kx7XonuLcUHhQmqPT30Ka5hJzD
yzQFPzoAGdgQ+me2Kklxa4u8sgrMNpcODaUQFXxKMyNgwZun/85vSJrbjo9x2L5G
MpR/bMMf4/cOIjy3bO4RPMD+3FX8oZp/fsShJc2XX8fL0/kCdD61booHmnJZWDpH
uAepsTPnvYsJkcYOvbMjLMEhN9kAj43/Xwd2Bn4Y5H+kKN2QzzqkzASkMtR7EuIZ
O/L9EDjtTbLrJduls+x9w/iJfOsc86b+JA5UabV5G5eDdsy9rub1wzAEKgYXyf7y
sY1Yz/7nocztSkNKHlTsZQoI7R/axvPMT/EkzM/fJeCxPrKQ0YBLrmAo/QXIMgKp
DeQs/ojXOb49XFC3Pu2fkcJL4CeY6Yrys7XiUxapQuDA/FdTSxUBZzjap25Bn+fI
i9Bi2bsUleNBM0MQPmVB1+pV9wAPFF4TWrqVMdIquNmQ5HA/m5CwxXpuCGqL+RK6
UhcylTTfgh0RUsMVTW9irzmHo44zsoUAkxy/zbQsvIePrGtN2yrSh1T++N/q1LSQ
DMH4p+qLTMEFkh8bArwu23bUHpvulJCoc7495ewSn9GuhtruAhg4lOoy2SjXqqjq
fslwV65MkTvwGoV95RvbGvqEnVvLBF9khMONB9MKbG17QQzyR8W70Yy9wFhVXT4C
6LxZzlRi/nL63vmuaxRDL2j75BN4O0AMm6DMAIWVVeGDof1OraiA+uoRPScJtfIP
RzCkhxH8KzSv1EFQS8misXyuPd3FuTFvA89K0TaYTcPVBEJ+OfxSQwwW7rOwIr4d
QDBZ6VrHV4rn/l/oVqy+av70IedlyMAZP02J0gtgMcj0mdkqS8mvmw3exTbONrsR
G8riEy2Dea7TuOqs3BwHJv0DuYpGEFxSwEkCKtvT8ezRZ7an4fejPDznyJIrEm7R
B8mfOz/t56UwNwJMr5ZjtWrRv2/oPZF2kvODZIeXk9ZbxcESUxWmhIOUPYJL9gBT
dYF0pVcQWqQMNlqY6AojfWQ4NWcvBZQz2tJ3rZfWEGaJ/yxZbPlEhDOrfYp6XnNf
7U9Aij5wGRL4mBOxPu2SLzEXcE3pYiU7eBJ47yaRC9aKpsepQdXhGp9KO4aUZDo4
HttxBI4Ub3P/EHOG3j/KSHhDJ5hI7Qe/Tyx25cn6/qd92lnL8g+mZNkOyUArU+Os
Dab7oBzCb7WaLKTW7Mm0qeHdMv3U0COF8cs8B00xjVw0DWAb7/jqxcxGF2SgC3zp
PEuGM6KG+GlpIv/FMCAiAtZwhTfqJvVFnw9LA8ZvgSikTDtqGxYkEVka0hECOt4N
OG0sH7wK6kM6Ep7wSLBmkvgLjoU0arvNX9/OBlxbmttZq/8VGIbAnCzs3Mt1T70m
TI6i9FdrI3ZRwYYMRXQCTUby05UwbvVEg/BjXCms3eUSB/bu8rg/G+cJFqlNygrT
elQZKJhqHBeu6Ff3wzlvQJUxJSDbludktrE2DwoFPltXUa/P7qwHmmpvoMI77p/V
+VtpwDw1pRLCa2jrdA8ePNE/usAYfohyyHeHYT7F5gx2x3AeOF4zeVF1Eot1Hd9e
IDFslkjuGox4AaCHu6ELKml+mLkaOauo+YUotnlwREH39Lz4KPWMW8etXO6IMhbf
xndI6n86hOpv94MRvowYiWWKFI+P0L72DCTeIdggAbiDFUqswbIamC+Mmclg1VKF
lAZRVkQuV7/qLILGcKle4Lxp7sle9mC88BiQbO9fPIYRIzPR8yLNQFNLPsLarM5y
gPuv1ihyrZmavYzJY0DlNJmVs9is7z7CJxqjnpnVfF1a8Z9XwCgAz4OqTK9/XueQ
2C+YsyJf4zbAB0klXXjz4FzQW3YME1HY7ygQtnWSBWZeUMFpOBuZpXvVVfEYDRt4
C3D6q0G5B9FinNl10q64ULdOw+TrXYS1+VmFQfbCLWpyMK8MIue3MzYlLGRIB0CN
YoC/APYn8s8NB97tAFFAj1TGM/JA5LIj68cYAXMaMKNWS8ckzzHc86E2Zy/MBK7l
yhn12vJfVDlZ51DNBbcinhDrCeDDhikopF1cHZBCPExFkKWFQbYP9xc+NEeI3O2+
K47TBmUMjTz6l6+4lwzIlWpFuYN4qMwoT8J06bV1SmzvE47euZ83l/cbJDeQMxcL
Qj7r5ksrDuc0NeiV64i4dehbRxp/ZMqKrJTmd0wbYCCCuqRBqZIJmFbBGK2aGyeJ
YCUZzovYNQ7jS+Q54EJr1TWewuOVANOrQDkxzDXBZfTzG/rMX9B4iRWw5yxNrHK5
Mrwz00XzhbPlOSqolN93x0iQrDzWgNeU0xoJHG1WSheF6qpAdPLyp05GHXJy9f9X
AbSQmDTDlZqpuzYbSkEHgZo5ZM7aNFEnAitwMwRkhLyBWYecVBSC9EgXeITB7Oj4
Qg6Ydhayo+ZuuB5AT984mphzlzIl5qY/RBZWfvC0O+V6f90uK0bXZplaDPkIOiXo
aD9YVLDlKiNy6gxSyN+HAPAxOb2V5vkUHOQwYhrgaLaxpQH/G5wXK4+DyPJ+Q5QY
cHP+xksrv92XrQZkph8MvUTT+RUreNQse32r/d07/twSPf0rcoRA8iTXcLqFPtWh
Ybp6/M9+73r+JuFKIldm+ntD5s2jZXhy945oyW01er2qznVkl2DbtaJL88s8yldA
d9q/D50RHdbhRKq6mzqrFfIxy7/DN7yOfdqclwabxjdjt7yVJgXaDDb/2pQURCw9
i7GnVT1ply2ui7ZYeGsg1Zkh6BQl9jeJCw6uHqpU128nLMS+eTu8bO2t1T53QCYL
rBVDOmb/EFJOIJw1xLvhmyCiFkkgmEqaV69wPmSCpo99tPXjI7NikJ9+MQU0SMv6
Z7NCmgV7ShSOyACJZX6mse5uKfZnnZAUxB/6kGyj7o6Jfrzpu5iwN3T6OgZjbeuX
IyEFZohu75txhn5dQ8O3zJ6Yv5oEGTCr/0vgSGQ7BjQKkLAre5HTj469sEH+zTBF
SSRj51i5P2B9hPDl6ksLrx8Ztgtb+vDNS1ETHaTiIwlpBkFFnhasaCWX0LerPM4f
IHmYrsXOs64SOI8bj5JMsl47V8jPdobuNxnHTAI9g4GrhsoT8VuTAnjnHMFbLwkV
n/vlIxnoX8zzxkmSfrgLv/WgK11aep0YAQ+cs62iAfiZ7xKQa83E7FuJ5h3Gtuhk
0rxk2ajJ1yyQ8o9sXJ7gduGjSF4CWt674SwRM5jEye0ZDyGJPOcyxch0tZw6VNo8
0BuMg3ha+Axy9Gm/sr4GLLMDQmf5G/IrXctm31EAiGLjICyA7dTxsU1hYwRbodgJ
xzvZQgHqCxgLyqw7BSkFuWIMLl3VJOgEXLYVSwz4fxrT64ILq/J79bsK7ocdwNlK
Y3TpR9PXpJjKlnUq0L8RDBREMi/l980/n08CUmyNj8AntFVjsIQmCNhIGcGpTWUq
+HZqWUZhAEZ3WncUElNYN9ZN1xD8usl7t7LHgwYofqJ9KJp+SP7pyTPPcFkgNZZq
pJXQvz/ggTiayiLwioxRRZ0IwokMJ941SQAUTemzvGyHtbarF71kD+45NjU51POo
KaWRayz0JIrwsIv9361S/XJgOq7pGkdEBnIert73sDszbh+GNBVoPzSaFSxN32xA
fYL5nodiENV99O9Rc2s+Z+pPgYCwldFxC71dDy9xMwWoyQHt8xcWyhpQQVIgiN2Z
PfmipJnjztxQpUy8aZCtIb8HZqU4ML+6M4mc0myE/WxFgnc3gzeH/8l/3yVz5Ld4
ItCKwTGLN6NiSheIqD7JswTA8X5GISo53Ts8grpX/3gVdoy0yfHPaK6dk6ySdeEQ
uWH9nxL4X2LzyntTKc3bszmqhqmEjvfI1VNg1UOQQUvRNkx2tNSzoKFsvFtFeief
NnN84Zyrg0zRlj0KOpJ78jEhgb1LyKZ8i7vJb0FphyU5sGtGfOPKQWecf9lQuFri
RB06Xf05yr/2lE/c7gwTi4dbiuWMRQ4ZEY7Rcj7o+gvapy5wtzJrMaMNQMeuRy3F
ERnhOyDK+uljlvQeTdhqtlp7Cvf92XChu4/hL6+XBjnL4NsP8drgzgwTxxrDpkJE
M20QER/kFGlNKMn+5fvFK7loNY44G5uSnrm/gXvurMRxhxJtgI+0ZinUKBHn2Qwp
cRtLN1cQxhcEsRpqzSvxm9CZnaaL/ghjfhnyfUTD3nfv8EqcvG4AX5/9E1AfETP2
Igy+HUGLm7JaTm5uSvT3XcPLPNupua+mF66skbKK6JlFDBCwgchH5h+7/79mrfMU
IRjRuCf+ucLNtwxo9jtvz2LGigtRyl5BLcOu0TP0/kyzJ2w1gGoQOv47PdzRZqR1
iSbxFU7wcpKnH0gxK4AgMUX3wuWPLyrrfFhED6GQs8MDbpyfXyMhJmSnC3yo02l8
/LdzDxjZ2tJursnJr6UmoDh1biNL9W6ssO+Aaluoko3YlfW7HQdgHuDUKizH+mOV
5baBKoMFdQunjxO/jXnAlUjHMhYiA/4qE7RYUZ88RcFbWBwf2a5sDyaN8H/Gh8va
lGygARvUjFQvtqkwxoWOQ8htcmIWrZU8zP4PRPCGsew0TWw0IxBxj0Oiskf4u34W
1tvwfqYFFOS0qeRTjEmBJeqOAN6ijv8KgXg8yQwOxGxyL8QREUPJAZy/cB7UMsUL
bIW83O9hTwJqZJ1SYlH9FVGlzxEoBvQXaQrXl5GtktWDdSDihKjbV3l95diJABbQ
C8MUdWBAJiiPYjDmPF4WmNbCc/KDnd5d7AsQy+dhGbTUlDn6TnDeTB8MkGXq/Mm7
Ovw7f2B/lZDEtMzrFLxyqTu7/pS2SOkN8TAvDxDeMYGBhW0/2UutX5viWhws6kIT
K6ftt9eu2pDqdnsFf1+FqEgDspk0ZR087bNbfJat+skVHn2bK0BwRVG4QxLK6nlI
jUt6DqYAP3dp7w8yFM3OP4dfOmhO68XC3rdcOTS3iFCDN5djrqPxqBHk+Jyqss0g
RnbACtwsv1bGqfxyYn255e0tOOaI/7j5ex7vR0Fx3odB12dfU7iLnwdVhP6lEaCI
knDxjHFgoocLSK3CRNWI2GvwHkr/MczNuPmeKHXqOv5voZ7kjK0VekA2v/WSOru3
k04+3LnlkHDs3Fa020dflv/J1pIVNdQsxJrvfwukjntHDx/qAK4Is10uIKPRZCHy
/kJD+rNn9gMzsq4CX7jGPHMviSgG5beGBv2jePxWbu4/De4QfXhTeJfQxbGH3VVD
Nrzk+i3K4XdEsvBuwgAtd1Sy9wqsys2jd5EFfEOXhWu7X6iPLRcHd33P+RpLYsph
SuTCNhzHlDdNJeFgQJLSf4jGGEpmD10H5Wb8m2v3wq/BFhMnwI+3OkZcFB2GD0TO
e41M4b5rKI69LAm+lrNCqNiEhaWc9nV5Vc2vMrzbud3k757rczikfhW/nOS76Q4d
XELDsY0pIX6qcEhQ4VfnnPbyIKrXx4Iniapv4o0VErJcBBMcauO2+BLG3Gz61xPv
KwKELwJxF7V1QFlbFi7+BCAlsr14pZVqV8QNwZbCW84w7hgaeCXEPIHPTpnn7jHu
FAD8unTV9A7SYOdRRRA49KAnn+6ef80OXx1aAQ3r5948jUa/HMzCXYTCXnYvkH2S
tmSm9dCpJVYFtjXuaYWEcBxG5RLcH0Yqv0sZ9rFrSarUKzVwghhESmQ6yxCSo7fv
HwZ9BuE4Cm0AiXH7lYqzB0YX0VKCQOAoR2tw7N0saE43i28yoeJYRtUEuNid9GoW
CiQxFINc6JsE8oH/o6MDUvJJHq7sro99ei0I8DbgeABNfbCVb5o1Z2q4EB7Aouba
yMhZhzEhTc7RPwppDSh3izLPHEdFGxYOp/oMIrPOlSqP5E0LjT8uSfnltmgLWJWx
70OfzMe4xF0k3mZqW6Tc6/eQroh98+pprKPtFRCD8D+aXRYLCKpRvuvZeYafXhAt
QTw+DJ4K8tAihYYU4iDa+FxXEYINjfnlzeYNkr+5Lm74rjvjc8F6OImYqTnN6twX
PE3hYYgbSEDXTVFmBgxnewE+deX3rv4FuwtxRDtQetDU19TFJLECVx7CkttFMxqm
y9tigicHCKg/gGJ7w9xaNUj4Ev/M9Ytu6gsoScX2aA1xqOMkMC0cpLPlYXL3aOiw
zgoLlPTY1w2OrfG7i/NilMWCl7/z4uQUzEZCgwMtURIkATHJS8y6b8KM6uQfqCxi
1S0EgwFpw4MIe8J2pZSU+noTY6vud8gy0jsuwICVBLPO8xNuJTsCQTWJJ4UuhlO1
bnxA1bgxeTW3lDaF854ByM5G91Zk91jDnriFY+5PuY6rgB+Yfng27HOR+edKzTqJ
kKrldTKVh3NP27KMCeY5+q3KY1g15TtkqpEfbaQnoZJ3DlUOSybyp7XMKzgUer1i
cZWfbgJ9QYhipzNVSaJRSh0x+77IBw+W08rJGIYPsgWEKdjivj8z6P6K/bUGBCOa
mgtlbgARK/jmSxspX1djNm2sForBqcjlOEm3nvDFkFz6fOnvrIWqCOP5hZloNGzQ
H/7wGgNAC2ciQFMSrNtei6ES+UDLBmfKpoFQtoZDTATTVMLUe4MIYzb7fw4nyGGp
m8WQcoHaP9j5Tk5CYB4LOS9SYpW/Yt4InrbMXZHO4b6GL/OvtqriEqjieiov4Tle
o7dxWNXrrZdMnmutj0nNOro/dh+vO6/KehNBjASp+BdF+3q0IxJp1f82XmKnr/7E
zDW9QdzD3n9doWfSjZuZsGd6SiqXHfpFBLN5oDwv3UsETrENR0TUkjbhcJl+bJ9b
1wVzJZwCl++J6+X0l+jTvUjZ6f7alBUhjy89FrfkwySTk1r6spicCftmvy0LsoVD
jQboLR28+M52gTztDxp/DwO8ZkorVBEpESudOG49/YyfJkH86RWWwBBiA/wmNxQ2
JUt9662B+usF0CDMoMr79jO1RpSbW9fBZ8JVuxoxtiHPt78TLqQFE4n9JlA1DK07
thOPLJGsb7otBTwy/Go8iFky7qLTaQD9lnIzmpWRt95G2Kac90Vs5kxG4AUTqhsu
9uhHdgn+OL8SSugYVWHYEVCmz70m1nuCySkH0Rvt2wJ+6K/zEZ9cdW0QX1ImF8ME
PDPNb2pGBHjRX5C1VHhIDp3z7RDm3KZLfg1QCh8xPf65tF2u/UcD2sWnx8VbGmt1
dw5oINX9RyZqUJpTi25GzCWYOb50u8MnokKTY27ZnZJ5E5yp6q61qItppkvKTACh
qKgMZNxeiZUH8cFfqYUVl5FOlidm9WfVyh4QuqA8eDUpq0ld6ta7sXiF/PINxThj
LPUXpWUGEz+5dPipzCSU9A4knR94c7YuAvHs2CUQJjOKeojO/sYi9YK+mlMOUNT0
ZDCxzoKUDv6zJinobjqSCTk1xRqZZOeYhUaDUfprFcGxKu6D2KEYH1LRG/+VH9wH
rTo5t0DqxwPZvTMOuwlO/sGpczML7hQOQD0xiuA3rio4pilXY2hKD5sbOtk/IWHJ
GBCByY2rLxg5q5yfl4JNs2E/pm+7mt9JuZahqeSVlHhk2n4t8dt2zQPh0zS/yaCx
LrrBy+xEoQW2Pi0nLPpI4DpbQZxIw5TE9JZtsNqPeJwHjNlwaIy2NsggipQkj4AT
rbWuXZkPBjGzgymL2x1hxCW7ZJIxv2WXoG3ZFxuMfoI1sjMnJuIgBJdLnHM4ClVm
IQrlSXn0FF5/ItJ3FmZhZvjD3GmdthDnUxAFML6nz3I=
`protect END_PROTECTED
