`ifndef __CNL_TB1_DEFS__
`define __CNL_TB1_DEFS__


`define cnl_tbX_generator       cnl_tb1_generator
`define cnl_tbX_driver          cnl_tb1_driver


`define tbX_genParams_t         tb2_genParams_tarams_t
`define tbX_testParams_t        tb2_testParams_t
`define tbX_drvParams_t         tb2_drvParams_t


`define tbX_genParams           tb2_genParams_tarams
`define tbX_testParams          tb2_testParams
`define tbX_drvParams           tb2_drvParams


`endif
