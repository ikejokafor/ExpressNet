,.mcal_rd_vref_value (
{

    mcal_rd_vref_value[62:56],
    mcal_rd_vref_value[55:49],
    mcal_rd_vref_value[48:42],
    mcal_rd_vref_value[41:35],
    mcal_rd_vref_value[34:28],
    mcal_rd_vref_value[27:21],
    mcal_rd_vref_value[20:14],
    mcal_rd_vref_value[13:7],
    mcal_rd_vref_value[6:0],
    7'b0,
    7'b0,
    7'b0
}
)

,.iob_pin (
{

ddr4_nc[0],
ddr4_dq[71],
ddr4_dq[70],
ddr4_dq[69],
ddr4_dq[68],
ddr4_dqs_c[8],
ddr4_dqs_t[8],
ddr4_dq[67],
ddr4_dq[66],
ddr4_dq[65],
ddr4_dq[64],
ddr4_nc[1],
ddr4_dm_dbi_n[8],
ddr4_nc[2],
ddr4_dq[63],
ddr4_dq[62],
ddr4_dq[61],
ddr4_dq[60],
ddr4_dqs_c[7],
ddr4_dqs_t[7],
ddr4_dq[59],
ddr4_dq[58],
ddr4_dq[57],
ddr4_dq[56],
ddr4_nc[3],
ddr4_dm_dbi_n[7],
ddr4_nc[4],
ddr4_dq[55],
ddr4_dq[54],
ddr4_dq[53],
ddr4_dq[52],
ddr4_dqs_c[6],
ddr4_dqs_t[6],
ddr4_dq[51],
ddr4_dq[50],
ddr4_dq[49],
ddr4_dq[48],
ddr4_nc[5],
ddr4_dm_dbi_n[6],
ddr4_nc[6],
ddr4_dq[47],
ddr4_dq[46],
ddr4_dq[45],
ddr4_dq[44],
ddr4_dqs_c[5],
ddr4_dqs_t[5],
ddr4_dq[43],
ddr4_dq[42],
ddr4_dq[41],
ddr4_dq[40],
ddr4_nc[7],
ddr4_dm_dbi_n[5],
ddr4_nc[8],
ddr4_dq[39],
ddr4_dq[38],
ddr4_dq[37],
ddr4_dq[36],
ddr4_dqs_c[4],
ddr4_dqs_t[4],
ddr4_dq[35],
ddr4_dq[34],
ddr4_dq[33],
ddr4_dq[32],
ddr4_nc[9],
ddr4_dm_dbi_n[4],
ddr4_nc[10],
ddr4_dq[31],
ddr4_dq[30],
ddr4_dq[29],
ddr4_dq[28],
ddr4_dqs_c[3],
ddr4_dqs_t[3],
ddr4_dq[27],
ddr4_dq[26],
ddr4_dq[25],
ddr4_dq[24],
ddr4_nc[11],
ddr4_dm_dbi_n[3],
ddr4_nc[12],
ddr4_dq[23],
ddr4_dq[22],
ddr4_dq[21],
ddr4_dq[20],
ddr4_dqs_c[2],
ddr4_dqs_t[2],
ddr4_dq[19],
ddr4_dq[18],
ddr4_dq[17],
ddr4_dq[16],
ddr4_nc[13],
ddr4_dm_dbi_n[2],
ddr4_nc[14],
ddr4_dq[15],
ddr4_dq[14],
ddr4_dq[13],
ddr4_dq[12],
ddr4_dqs_c[1],
ddr4_dqs_t[1],
ddr4_dq[11],
ddr4_dq[10],
ddr4_dq[9],
ddr4_dq[8],
ddr4_nc[15],
ddr4_dm_dbi_n[1],
ddr4_nc[16],
ddr4_dq[7],
ddr4_dq[6],
ddr4_dq[5],
ddr4_dq[4],
ddr4_dqs_c[0],
ddr4_dqs_t[0],
ddr4_dq[3],
ddr4_dq[2],
ddr4_dq[1],
ddr4_dq[0],
ddr4_nc[17],
ddr4_dm_dbi_n[0],
ddr4_nc[18],
ddr4_nc[19],
ddr4_nc[20],
ddr4_nc[21],
ddr4_nc[22],
ddr4_nc[23],
ddr4_nc[24],
ddr4_nc[25],
ddr4_nc[26],
ddr4_act_n,
ddr4_odt[0],
ddr4_cke[0],
ddr4_cs_n[0],
ddr4_bg[1],
ddr4_bg[0],
ddr4_ba[1],
ddr4_nc[27],
ddr4_nc[28],
ddr4_ba[0],
ddr4_adr[16],
ddr4_adr[15],
ddr4_adr[14],
ddr4_adr[13],
ddr4_adr[12],
ddr4_adr[11],
ddr4_adr[10],
ddr4_nc[29],
ddr4_adr[9],
ddr4_adr[8],
ddr4_adr[7],
ddr4_adr[6],
ddr4_ck_c[0],
ddr4_ck_t[0],
ddr4_adr[5],
ddr4_adr[4],
ddr4_adr[3],
ddr4_adr[2],
ddr4_adr[1],
ddr4_adr[0]
}
)


