`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sAe6crON2XHziwEvRRYZF6rGps8k30he5vRZswqx4PODeCnx9QF687/TbRWDKjXE
ZccZPrAhh6LaFQ8tRC0pKQAT6cZ5v0VTgfOHziQyKSyv+6SgiWZk7U34OOYgK+Fg
r41FYLGQM8JXmibc+igGEXq9QwdI99f3o+fiG6/br2C6tMmu8O4pHGhnMzb/ZXYX
RfH2dSkiHfi8pihDEk/V9ad3jGc31F4M+K9cZlqg5J2ng9Xj5F5aEfrkvhr3ECH1
Kat3lZl3htkiKZBLpXzdIDAuoryHtGK36ppR1bSb4YO1zmnwCsh/L9F5xfP5crPl
clDU1n5PfyJPPoB3yWF67gH08qXoTea+F4HhF4e1UQKN5qJheELjcZZQ6thPGglm
PLOLngeP492oyBINxbYEhV052GHKDYn8g8pNA+iX4wmUd/3oTkpZwdW1gKWONiKz
TqN/d+hTqB5R/CpRPNXY8iuUJ1LE5CoMD+TuBVOMDl7QOy/AoAzKj/j8f2qNN+eu
tsbmwnWAC9xMeJNspZZqRB7Go8JcsBxQU2E4i/CX2aj1EFyFgpK4HwUTuBzy2p2R
bMkgpTHzl6kvxKOCTwIkeceHfEr8kFWWHaaovk+Du/zpCzJMNxjw7K7HvP+Wsi8/
OERsaUq0xWuMh1Cw+VT0c9X6a/A3axBk73XOG2fjchWT5xy/UELOep0SWGj5owkB
r/+cNBv9NW5PjMS/R6K0lH0R695jtZh8krx4o3Q/rgY/vFNcgi8w16/h23iAdtnx
Iq1CvYZ097p15mLGjuf1iSYy9FSRntfHInkGIdEk6qGobS9AhNjOz/I0XT6j6DPT
IL3+iucLw5XXDVGxbbghvd6HhTCYFjGyu4TzTcTE1u8X4lrLHLFoRA894Mo5K9wf
k0bkxJreONWETE3iGUUXkztpu0X2LRMBmt/3kYNPIjZ8UhNE7NfIr0x8EBQCJJ3C
XtSZY4BJEuvs/2pEKwKNpSRA7NjcoP1wAgILWhMnjAMmN8F1YbQS0gJDk/fufnPo
t3UynKDgqzj5O2BIyNigin9wQg26aAQLgh6wDbH5U6kZll0fOvaNR/wTx/FtMZ1s
2MUAdb+Fy1Du+0kIL8qpqfVnJM7jhHQq21RZv+SKed1Lsrsh7r72vxWZxD7PIHkf
m9MXFIKt4bnF6b2bKBiETJkqdkzrObo2hsn+srP4m/xlEw083gNV48DdnJS7Tcx7
QpO7lFi13rEwWVqzT88PnhYCi0VY2119q/aEyJwdxxL20LG1EigRhoC2P6l6PyCu
BPKolSty7ZP9j96TnpRePZVSBgeddfAaC5Q6aK0uDdU2Krw1Upcd/GEfyv4DFM2L
JEtjMWPIVqMZDF0ZuaU6KwI6wpAoW8bvTfjDliuom+fbZ8GSDcD0hx9J7Ifnx+xq
KJmv1M6k8yhHQcz6r32I9oQFMS/gkz5VRA5/ZIkPoS/h9+xEf8bu3+56lqQABzst
idrhXJLuAEy6V5KYPWFC0NqvsqlGd0yh47dxmnXkrtbH71MDVuDK1Cw9jtXQuKvK
wqXDd0YWhM8IVhGP00wJtBY3F1ac0qs5sAFoA5G09jMjI+1SESBeKLVy/d7/NEVP
GRIsRwa4TxlgqJ4c7NT5KBT49dFYwe77PgWFA5iXG+gT+G5IVMilLt+skIQt+5Xo
xmfpvOpWqdlx3sSyY+9kizf5fdA7blCBXixK3yy2JwUEGPRe6ndCt/Awi6wx129T
+SMPsCO0UQomAzi0YRIFN6Byia5ct+uWqbCRju/PDXbK/tj6otEOWvdpZkNYS9PW
WvARn8z1AtYXP1NszLMIBVeF1tHzO9ciWQOTSEWQ8FcyJ+r75ujH1eB12SIvoA13
1KEtRosQKUkNv31UNkFufRE4zLzJp/77TgHCXW4QHoWH7wmJjOPqKe5eb++eMoju
j7ElE2gM+/RX2naC5B3Zz04Ipeg9QBGFTWI0JWNFw/PFN5v0Gd1LaGkqDrA9mC0r
nb06maEBconms57PlTThHGRl8ZKau5DMpDiDjC3m71V8hsD/WwgchXgDBMa2n/9C
oZ2FIGnxHIIF9Wk8oSP5XGjsM4OQas71NTknPgiKYglDCCEtSgvTZyParO37nmyP
Vgx6S1dPdvxFFnN83aVpU4qj9OGNnqaTWT0tgIFAHrD2LTS4LtexNk45ePWdw7iT
nSnRi1nl+lgamNYCUUg/gi9N6eekIM9++8XlYHKGEUoJMc95aQaRr6jH/PQYBT/P
+ber2BkJtNAesKnAgz0tsU5cx0IpYkkq+M1o5D8vM6ZIcBBONdOCmUWGcKhk6Tv+
sQ2p85W0JF/w3+kUcNal2efXRABcjJ54M24TbKvhBiy8k+Y9ShRIDMqdNFWJ13O/
dcbi67RJ4/NowGRS8U3ex8yHQffX5+2FEgTTNgwrOLnmgGkzvhrxIC7XyWa+tON/
YxuxMyTgfQRGs/59f8XORAgL2d93arpW1D7QtAN3DWy/8p6o+0NiBqbRGx3NUJam
avggrzFlL93GUqZVCIb8XtLhIu6ok+aFY4VhqdFV+9niuUW6lmOYW4a+1zfE9GWV
AREw0FKXCjWz+D86AQzrbV/qR3WHDK62nCCc0o8cStOyekGQm4cZ7OnuRehY9Ryj
S4SEioMp0ai3BK8EtFuZNGAZ/G9/dTs9LReFoZ2s7nNAZs1Q2nvwlKTtnQkaVUzp
HFUZEDvUDgU9HFbdPpWGP/oiSAStWH0i/Uv3HxYW7mPVVpg4ZgB0+mCnvPCniaDd
/pzzEL7LUF8FvtJx7qZobv8KIAp+N7bo2DNszhl/1KHxJIL0zIn3M/svSLZjfh/f
s95mF6Z0mXypmiiVAb9M/LVrAk5rbmYJ8QNTsxPJhqYfWr3pryw6fSAImaPU8ElH
JGhq2ha26IkAwSu2xfdyxYKzOUEiwdmLDhT08THZSd14cRsaXWscUrKvtqGXvJ6G
uyH9bPn4shJYw8qw4EeEaZXdoxF3UxE6ly1DsF5eu4fh5b999RPetqfRnmT/G5MW
xrDE+S2Dki8wFGx+P0eGkT+YY0MJYg05gwWE0lADp3J/zqs2yLDMmNAspoOC6F8A
k7syuMsrU1I0DpnS7CJZ/UAD8lDEFjAaMq25myxra9WvYhUXQ9j+hq32utnmx1Kp
gLwDIDEsoTF1tAcZ+8GpbZuXMlDBAHnaw03HTpU+i1T8DVHB5J/trZATqU0Mdrw9
h+k0F90sZxq23vGZ6eEboTFhM8Wjovox+fRux/f6TbLUoyS6KU0nAx9iCvcwgCzY
v+U4uLTBk9346BaycdDlsvpke28ynIa9F5kRzeePXnv4Zl9n1H56eqgJn5VnsRcl
PD4h5ridcdGVOYr0fKSsvvws2T+9c3GnYLAMG2Q+JC3vE+YZvVJEV+3UDPXQzPh8
P9O/U2SStHHFo1JYw2DAGRq+AV89Mlf8PlHzVDX9GgChUFPPgqK0Q4YfGipwh47k
6JMiC8aejcZc5YPRUFlByQ+GAkr5zjrBrgMeOuX340tk3otsZvS3p1JN01fye+o3
K42pzAszUoeJSv/QU4aHp9XxEPzEZBsCBA2cF10lvzV57UfOQpnNSKcCWcyIP7+t
FBT0eprfrCSFY4AkNsyZXh0zXgOuoQXouZYeE8WaQ1HKW59TorpKkRz3N6Oqe1mM
4w/uCGsNMX3bOdrE4J3S8+cJlvt1pm48T2P7C9VJc7K0tm84/T587IE14XCIw5u4
/+suEPU47g0tswCa+lC0zj4//KNPqQFhxuzSyFCJJp2FmMPoE2vypJtGVRPT+CiR
yuwLfZpr113YCTTAiFWmfHGHGL9UjWV0k7F/mUbQQMwrPZmDUIM9HSe7BHf//Bmn
HerUrHi5iOACYtTGMcME5dKkSshl9rQwWql1kOZ/qJiy8f6+E4/dXtqRSwrAJsVu
yPLekXsaEbu7J6CP+L3GypEABjn93ekH01DWa4MR92rUDxiICfZ3HP9nH0soxmVY
gbXISoQtPuuaU4OY36ZCF46AaDmtUxOgLcmX8Ry9uC47BuU361NCxVc+U+TYcGfC
D+LQKaFjHWYTkz/MZbCPPQrrXdRpFUvga16TNlPNcG7oL+SKhm6i9XGFs2Sss+h5
CHqXkbYxAMNrHMXSqAucSEMQHg/qho1788jEqDF+g7OWOxvUgLY3IYE7D0FkCTuM
xctANAcpSVZug21s6bQhVHT9BRR0RDFE88/AWYAtBsbWFyWwYc/szLn4wBoCZAdy
vpjBkznUL0by5lYoJaLqpFYvfOEp2ekp6cOJIzoyD3yqDV30Fj+ysQmKce52B6YK
CmzYf61iewhAe8ZxVs5Z0zFQ9+64SiYGxi4JYuuwE4vgfX2lBTD5GH0ol0nDqKbv
6XW3+6ouEe/FCZOJ8Rht9X5iE8qRNeHNjdis3hlCh1amkdnVT34+XaybYuXjpb4A
FSwQvoJx70qcCZLdx1SbesY5gnPj13J5l1S+76GHPgPGTGpmllHgepC/5qvOniO2
S2iYv4VNosDQ1nTwVuOeKmQYKcHDV2hT2xLq46F8WJfeY60iRELkwcePYVA0Bf70
TAtNm+oZFaw4dGltj16JYxTUfdNr5BTfl/RLOcQX6O3nNxMqqf4D2PZyEJDkEdqR
ahU3kP5yTBGM2gKkBVusJDs7t3uNpmAvFCflgn4yGR0x8/VJEIDIRbCXNMvjfrgg
Fh5dR1kpYxqTMWfV8m1t+YyOEgj5ynDM0LohDcOExD3XpHkAk3uBApLqsdo5aokn
thZyQfw5j7nlJiFsXhfFoZqlk4qP2fRRyiZFvA42yk8xXqdf9YkBHwPRUOsWT55m
/m655OHw/Obaxhagz517BOJ4TQzSOaG22dt05d1PJTxbPo577TunSuFakI1MS+6+
o3gtcne3KrvmcyT3h2qGW0rAEXTtiq7weT3JHoTDGhTFDmDciurHIwX02rekiQQy
RQvUKBOjO7Vz4PiwIE/Ls6vY+Ts77BBYo+gp1Faxwy8gZ4YRHzMOe9fu0UoxM2qc
BYsF31rXe/PxquprqlMrzvj/ra7GUVDd/uFxrB5kgLzh7+e+b3AmF1Tm9/IkHC1D
qW7fd8gsn7fymHJdmwMXB2hkSwtW7ncUySnJN6UW1vI3tqrOhEkr8DnnOEFw89AA
y56SuJg1qU9QnLc/cTgBzkyGqD0OJkft7LC0kPqAw+Hr9A6wpiXiXGbN+mdco/5z
gykqu2y+PNwM0yOmi825iJSMUSyie8HdvrLtkjzjW5NYClfC3yV31F2Vzr8k0zd4
qslvv3PS9kO6zKKeKQH7PWGSxotgcgYHZZQ64PVEHpzQXP3qsfA8IPRYDmSKCIAm
/WA/ZhTDZNpC9DAsbAmq7SUFELKhyJtLmHZv83AaxH4Zv8Hfax2zolWhsYJ0DS5p
HSvV3R6xuLVYohPvASAlf6EMD0FBToISPDIT9eTnUoynTmVKnuDxCq0thPjzYnDQ
iAz20b3xJ9QQ3i+XQM5NgqSDIBQqR6/gRPkR05x6pBHVKlXeVNXyxVtGAPzoMXZG
BBqf4yH2xdkNSzUvXPctgiGzUktPAeSRWCGCbFkRdkARkF9iRHgmtxUVIF9kqKMZ
G727lWb8bDEtRQPSJkGJYl45/o8jO+Newl9qsuXC8PulaAmelAm5mvt8q8BdUR9d
AkH8f9vCgPH6HRllNpXLbwDAqRGT935DYFhwSF9jW9FdLxv13vbfhM+ZrgS5l30u
A76bYv9R8NUy6RR5Alzx2FD92zTYXzgnUhQ31aCGV3hbWWH8hGt9OzYMMWdw7RIN
fJBIwSlijs4DNGN8bcIeVzm8HZLZpcRSphl9MkuWYVREuscJc4hE7+5RxENxO9cQ
jSAb9oXmAA9XFt20ALVieC5Q6Wpws4Nzb64BV24NIQt4H0D7mHXxUBTuKuOamFg7
jLholp1VvQoG8kmpNrlEdtWaD4Z1iB8ETO0MW2buSf3y9WMq3m4qRqAb4NnzLyi/
bJauyKyLi6w5jiU1y6JfIi42FumV7uhLI7wTxUexVgZqVKFIIv6+Nh7hJ2cb+cWo
jA9PlUzWlaJecXQYSgFPMQ/EtosDVbiutbaQS5lDmnZtfRxXo79Qv2A9LhuddPqH
QwSm31eWst0XyDWen0hDPnWqZvWzLBJtPXoIJprVYoxHYL+3OR6lf3uI2o/PaYTR
EQKHSegqcxzZDCaF2/mFTHuOwb11kdBYhgcSnBIOOySlbK8L/qFQKhOTcByMNp9F
l9UWBJ1z97Zu1qgcQmDNpi3zJyV6KY/Ppb5c+GXAfuPq8Cr7Dsa3jdU9Gk8h64vj
1sdKLOQfXerT1fFn2Z0M46QPP4vO27r4agD6APi17dqsia4VeZmyJWh880j9dQN5
m4fSPAGP5X2gyWo16nwK5ze7iC6SA2EoA2vPRg+JrJZo5NiQorROVTk9E2WkETVQ
d7njnFYcpdR3X8VvPHWp7khkg+yoD08mQb09cxA8UGH9Q/6iFn+nOPygN95/ypjx
MOlzNZcrWqz6cc1mCAHHXa5doFw40U3SMu6B5fwIGj7olvLwp7O2pzBLBOq6NfNu
qrsNw+/ratiTMkkqGYXPPmRt/sCRLmmeSxCYf8+BD9j5OHT/NJXLCxZyEa0UObLp
sAhzpU87XXUPu8JTQs6+GUd8qv3BAyPI2ndPPY1YTA0BfnUVODt+GhteiUF5cvmu
ZGv52kXNf9Y2RakIDcSCzhjd7POpxPBRRR94yVLeYOpliJ0NdehSL+e3qq9xh2c+
jC+mF2EREmg5mdLu6O8uPmECl557QGLa1lV4Yj+kMRhSA5roxp8Rgi2iIBxdmgPC
s/rytJTHUIh5AU9s/orpplGv2E9EJdAR7dnQMn8qnD64dwbmkylssQfzepD3Nyeg
XXcit/uiYKZmDPSovTNKiSUHJ/fM2gebz79xSEO5tUe8SaMMpVbhpBblC7fwcR9n
mPMFYcQW4uNap6lQj5r/BeIwjeX2ZrYenqrS4CX/inKLkF65kq6qJ+2rn4X8sXze
q9x3362q2KBVuHZQJgkAbfvBVzQgFSYKePa6+hJazMPDWzA3e2Bvlor6EL6HTHes
UI9ovxBKzhLIwSqzPD4bgRuVPNdD3U10587Fu3JWQ4zMXgYEwKblkVo14HThwh+I
obqBHQROb6dP8/Kf/YQ5YiVTNRmZbWLHIcDPlGr5HfHLgaOWrbBgRCTDS2GbA4gM
6GOB76Ov9z+lfbvxZQncoPGAZ3RmHrySvAaCRrmHgB38iXN5aYBuigVZIhLyvlES
6/3B9OZRkei/3DH0Zfk3jTSxC/ZSBm8UFvrMLduA+RTvvidq7kbiPFUJvL2O/7uC
OfmpYzhs368dU3nQWyuQJGpgMw2cv2KmJLLtO0smJLgmp8zxOOmCRhdmXSqHIGIm
0cbKuFovXnSO1VR0QGNHSw2Z3Ulmq7iGOy7b6C0RdMMsD569avHd5sAvbBTMldFM
hc5EOUUyGL9fLGwgEk61mL2sSuamwhdtL8qjCwRrGNmnJVtxVTA0tjwyPPaXGMDh
71a99xUOYPCqfoEp7mqoGXXePxyWup77fF6HXLfP6lU/mhQ55H30h5AfbZ1cEMzG
T0UPSsZzdEMCzSxgN0GDW3C5BYj5UpTnMT+aWgTxLMBflpQRtzCmYWQnfyEz+ux6
BJVn1/w6l9k1+dBST0SrZP3TLK2ZP9WrtKyzPfFaMqFJZm/nA2K5m/wv1y5zT0Qw
MeJeD6rNf6mvNVlfESzWU7Ml8Y74SVsLOlf//JZYcqPEowVv78nDMQKDQ1Hnnamn
O26dECI5hEAVpoU+j0BWLijPpEFgeAkPblUluBN2MbszmO6fJ5KRS8QaHz73Ewz0
zUBIF3YnfrMBLZHyuXS+3nznYMHfDcWA1uEBbd3BxqQ9QDIWD6vBfOztmhfIiZZl
QCCRNx3WNYtFx5941uNitMqkFsKyCTrREvdywykZCv6Qk7PVvW46IUr2CX0NObOy
+G+2jPq7sHFusLYATuTYFXkBVbbrnu4F2t2Fra9NWeoaGxsF7NGDUd07vvsFN3if
/HPV7r0vQXgG6ovLD3VNcpuehHA/S2jXI4LMbVrtmoODb0whjStZnRp6mivh3+LB
juloy4TC0kJFCD35Yr/rH8CsPF6zF2OGQj+U8UGl8dcxkbr3zBJaFj32tW6/LyLa
airCTuZ1j7owhkLkxgPu8vRf3FG7AspVDvaS3cjXobkw9eTPUTHxutJml8kOhSJw
P7ekkn5s53hlG9FnLekWhStnnmb+sY5Q1zGPwmnAc3+eKlZXb84kvhlaGSokuA0b
/H48GOOd/65iEtuJ9llsW9NVpxlXTYVmWoH4DQ0CgICXHoOtqT04RfNPHGdpcqlN
EMRqKY7w+O1q9wbFmy3/UHt16X957wmQnWP+qUSRSTZS4GLjanqTxJjq0E+mtF14
X+mrxpkiXgjGvi6udJv9YesgJlnRg+6rCsi1iJ8akMhWj8nboRlfnX+JVKCgxEJH
dLq1C/N+L5CzdoAOSV3S12BBzqWYXZFxZk3Br2jcYxHWqHGi7sXQKW4Uoi+WJAbH
vWFJJ1lIHcfjhTFNL1069nZoe73fcnfY6w6zUW9lxFPnOWAEPO019E/Ghh89vjpn
7/D1/WlRd+gP34lWhYhlR4/rEed1RgOW6WDFVwsBOL4dMPoridfLoD+kcyc3dO2e
pn9gOYRmxyAb2I8BriONyI1KF5EoJ92/tOuezVam6EqLXb7uc6I9RCXkDXJooqHM
aqTzW5ffGyjZq52e276BbvBcSPH2KwlNa48t0VztPHeeP7YjmFyQcWqTG286lj0g
q7NOWg1k1QLgOdW3cFwnZFuJ8Ow5gdC4UfxALfvygNDLCc4NRfbx/fKTTq991s9K
9Ltdqu+Cfz3FdbInIqm9TESeIQGFGyqZjfb6JH/5uhxhec82xacW9WntVPYWDvcR
/j1CpsRaNtuD704uN65xhXg8wWJkNcz/tcBM0PThYTr4dIbePJri9TPaZwDavTlo
upKcatyARsHMuN9eKf31eQRsZBUYwnJmaG+Qe+ykHeBe84GVxxBhSemVDcRIPsHr
5a1VUR4kxfV7ce2LscBkexPt7NWkYpdh8fTpayZaZxOXwhZMKpalj2Ggpob6AaOY
lCW+bQ+AkMP/Xh1r10b0VlIh23ZLYgk49eF6P0ouvYUAUR4M5DCY0dTFTboyoBge
g5sDSp6fJW93HWSYlmw8afoaQ9+s+DgQI6FtxOVi1qNsK0CpGZlICj0TooQQ+3wN
IRD+v7thViIfmy4sHNaGNXoh4dIskOctfPW7qADb3qaB1Cm5ah38Dbg5OjOds6lf
eyfBTAvJC+Pnyhb9jFDnpntLoWblqD1e178SquApuC9UWgIVfeBy81cixsWZuW15
thWu8Cw2YAyNmbT9BVVkoudXsMSGnfDWt9qpwoqngEhyyeTEt5dddL+82QnkYsWB
RP/rIdVW+ps35EMYpVsNmM5p4xYYCgUmSOU0UqxXrsWx0mfnz2dX0uJeQ3PWvcih
D1LzDGF9nBUaz5J9/AYevwiLdBuvmybyRd3Vk44/onYKZeAZNOoW5AXTKSwIlCBF
Hw7devHUmNZ68zXgtuzP0eaBG3DxeUHazlPq4D3CXtuxG2FJC5Sayp0snvVokznL
74D54ueJvvNv3PkdTB5TrP1vfYkOblvGFiQxaC8EINw6aNnmXWl+Of2ME4m7jt1E
xVgZhnJcKvft30SdIbnfZ/6rnj7CbN5eMx+4u2bITjfS+7l3Jl7cKwYxyk9IJTvi
X4JxbcasNZag9ZDy9+5KRlUz0nO9yJN82KZeKEos65W32UJkJeLliEtt2ZKeHisB
ZkrNYBSqD+km+76j/u5/OoUlyRdw7FxroW3rbmgFnvxIgLQt64ibbj01V7eIZMWN
9ayvH9UsJ6eKFfvFERjXqMNGJ5BzU5hLyE2G4aS5hjziiPkm/ITL3O+e6yEczEVm
wSX+wqt43lZVYxGotyes3POVzkBKA8/AyTu5Oo0v+M9pKL3m3PjyusHoJZEm02Cf
cCgkSjLMT1NB8jqCX0JHDFvPEU0QNqK6hLzGjYJB4dFzZ+iOpxgVWZ5Oo7haxMBg
/YmlBurQ4FOK0y/P6rIMneZNWOETmT46nYqyHPGkwh1uGn4F/KW6f4TcktXQRhpZ
k26kRqYy0mT3cPf1zpy8gcosXNnNprkqjMZvtHPKS8npo80xG+8lvcSrdwA0Khrw
wcMWwpi6zxfIP2X0R5QZA5w6afJjx6E/o1phRbOr5KekQMNKBy9wtkR6IhSkhv/G
dFpEz7U6O0RyB46aMd9ffvGZNO6Ahs9701QU43ULxNIgflmuWDDuTjDh8HJn9ABf
06dJ2BRoRImtzNHwLQ3fhmvKn5GPWkTrVJqGerraVI0zBmYB0VuXdcLTu4EGfeRM
/WQ9EIV8zKg68gb2y/CGxnSrkcXGYV5vm/+DX4L3dSOZUzyl8oAuB/Y59hqmNUx4
2V3n/zKCtg/tbnQr3uvl4pnciltOik+/iYcNTbFWKn+T500+AoouXtd4fas6AZ+M
G/UdzSbM7vyTdLYhitQ+m3dMQQfG6ttragKri9IIw70/bjHdLzSz66aJZUQgL6lE
rY8D0nvQ5DucbscQceJ1+q1UXOS6SEf+zfFan3LiHArumeEbhjhgwCr5PQjR7X2N
nCEeL6cNq1eMrXtMdEE5q+KyeGb1FDqXzKOXF91ISIE/oHQZe1cC8ypdRi6Hz5t5
+uibYhQznc+7FgaSo2SfcXQKPlv+5k5cLj6uZK/xkTx9WXizfUlPpIEIDjobLSr8
IuvQz5cEcVWIv3Po28EjFpJ0A0Ha8imKDT+2JY/gl8/qD4U1F45TSIc4v40hYtWT
Ec01aszpwqnCJSTt63DxxucwjV/G95HXbSx1PHDCQFoAldKFu1tR6FuQsbh2PfDm
uFHF+4vubF7ul8xLMSM8LqehV/Zw8IyezyPLQUTDSbQkoyEHg8i0zY5xd7a61sls
t7IpFAGBIpC0rq043xq8g8BxgqM16d+fGlavpzS/C18ARN1nwepz/o2wUTCmtnAX
p52Ipxh79kyKZ0TR+9tEz7U1K91GaF8RFGlrlqerKetyI6MrY38HAza+P6STAf7O
hyilIE8iiO3fy78lKuYHhSjDKyXGyfredk6NdY7BAcxtTomfVocP/KOVCUgJP1EV
eW4wvm7JfONSh3jN1zXFCT0YfMZ64gWB4F65/9T7BVeHrrYhq7v2fp93kqAzl8+e
AMWYL74IcpyCf8gMAVSc2OAtrXAwxI3yhMmW5HMbZ7Ej8MDDuaQL00NEkMjDSqcf
xpsCNu3QyzyY8+kG+oy5QMQOEQ8WLOoFtlTiz5D8MsCJZEY1JpMY62JmLrARNsVl
GZ6xp9sNPgcstDVHeOimmSNaufCpaLNu8dU37ynZwynnDNlWd1mZsyKohOJLwps/
OQJ9VoyTjCZASXyFJ8rd7636NmUpZvgiEJSCSIAfZJ0mY6gJG/eSSeg+EXUVsbF/
AQ4kZ/cSqd+tmrd1uukzQdzdPLpaUXW89U9AQ8WNiDWzgbsQtEDxuPya+7ixGr6x
jBLjGE+CyXPb68+oEa4Bf9Oec6w4Rjj5vSpGUO4z93uYjnZ/zsNOfymm1hRfZTZY
B8Y5MGEij9B6ObY+0mq5b+1pMNBvhVM2KiDnm04KaZ3PNNKtvVXVamljNt/Od0Z2
vsn4Ej52hECbDOfoDIooVxglnCz9nMTakppKnj6i0kz8xgdOdjzUmDmPA7G3rOTg
BZDIXCxEGevaDdDfwmVJME0nEOtGrrw0XwPTrXmlSJyWrEPmqaJ2wc1wSEHI45Bh
OD0MR/5/InD95LbJy3kYlm3C+We59KtbBgX4dBbIq/2n1ZE6ufwyZiqxXrQ9KqY2
RvateEZa5nM0/xE7NgntNaznrvelO5c4CPSasTylxhe9DUquct02fCoNCY5HM4nq
TaYMzNfWx/cqEbJS+GJ5+Y0QXfioU1uvM+Ft4/rMBQ95DNL8kgTCJrRNKxecAPe0
GwReMcWltfV0jhVpytbvCOi9G8qWEZy2PHC9yKxwE17lHt47Fs8CxySHeqZ+6wlp
69j5/wqvqxyXC3VcJ/4iHgczZLkHuYnK0wGdZr5UEli9V9bxdsYddcKdzcKXhlpb
fn8QMiUV/5ONFQ20BtIQ+F3EzGwLKv0pTPjoFe07UnS+nrF6QrQcBKPeidAI9hPP
s7euRmjzlhUIKD+xGMg6b5TTPFz+QfoKwoXb99lF54vYqthYnoKMrzzjV4SX5fG0
+sLwj0FpLJN2TF04eCesVhdvOBqG50HwNGnk2Rip1X/CqAARGWGCTPFrnD2LVDQw
1TE0+3b2EGV+WIAwj6kDHKVHSWAKsLmXpOU7RwU4hVrPVmCIsvvgilRzlBJ3UKIe
IfAqATeVCS2OhlT0Wvp4e7H84GPvRp+Jixxnr8bzR0SlR+7OSdlNd0SB9jf/aXBD
ciHKoe6l100r06cpIGIbYZKNfIKDSPisdYLCmZqyUp4bAvjXGL9VargeZezx9/ZT
SIPts0JbZlbwZcIbrlTM+8lEJtInqV0N3wXXF8MZEXqiSSCYUIreThZVu11SFbIB
jsH9Us+W/MfB71Y3uCj8co/dmOUVZ7yCHuJq0G8HrAN1O3mKcVvas9fwo9rqs3eQ
RPUK3ryws4Eo7fZOGaFB7UzzBlZHWU0ZEyiwcBQdHBit+fkijwYSLoijWHeQ1C6S
8bZ8eKOKCyN+SHWpNErR+IRxjWfEjdLyFm9blJrJLO4YD/T7P7Ktodc9tP3f/xJy
r0Tm2Ck9IWnyp7wm6aBAqg1nas62EiOM9M0aPJWL8YxBCDITfDTTLkTxpRg44f1E
DOIz2r0xF/LUdV3l6LN4bAdbvbQPa27CG2fAIUD0n5hkkUD3+Vop4RjIWVpZpjSj
bWKlmeJnHQxUtV0Dy2cqbV0PD58IJHTo2Q/xTHnAHQdWx/JTXCByRwkukUbbKPOI
+V117MU5cAH/bhXBahCulzkbcTPv9cVvYLh7jlOrqjW99xxOXKHIwKocTfAygV6E
YOtqa79nww+zypHEade2Y2cFTwau85EukwsU/uJGwG4OZU5K32DxlXSgR+1XmNtb
LiOLszx29mUHVuOnH4s898vMlXRBJM2sqqr8778vX+e/A+HQ/Q91/bmTGH5btIrH
A544L5mzl/aguOzoSfgMOqX+2pQMe01gL9kFzttVfvzHBqrm3bj2IQoLVxDZfiVb
RxrW4A7VGvFE/C7iug2MtsPfJ+mz0QZuYtDlqumni1jjqQUyiCEdiYbUMqDUcqok
/X7L15T2rlCN/icwLvzP07ISgA7R/aT30xUNB+kHgylOjq6drQgyWJmILYiGmdxF
w2OIRlyUfk2ioK4WveHOJT4WYneab4oImj6Fazo33SZ5VcZxx/iEVYm8v6mjMC2t
+ahxndEBlD3PtLkvo0zftWbEuo9pnycxNSbmdRL7Z5I0dHsWhAQvkQ8v1FOswJjq
ilxyrhh6Doo7Ix3ai2ZQK4Qc1wJP4/Qcm+W+Tw5gCOOqv0pJtpSYuBzaa3tNNWBl
jnK+FAgsqQbfcHJKTJUMQfL/yqV7CQd26rwUEbtJNLgII2bLNcezWDSaTy4w5MPq
Am+yBWCTnOFoZHV0DEvIvRplLZ3HUmPrTpsiGkfc+aD6ySSsGfD3Z4rZHJf5+t6d
XLVGRxstapMEZnQF3/xIxVtC/CpoJQuwaPTk/RyubHWUhNy1aHslRQalQvp1WmpX
Ulx3rvXS/bwUkXsDAu2RMM6nZlRRPLGFMCYhDnyjmDi5qGb6Idz6A9gzLs8nlVNV
Imv5dyX+mJ63sriUkbprdUG01ZisZ5G+yIX8joOfi/YXOHMFekH0O/bu9HHDj/pR
8bS6K7XuRkTM4ZWMRLlJdd2wjDXbt12qh3P1mrAguie1kpToAHU0SkyK0o/6Jxdk
F88/RFzslyiJfa4XkBV0WgRGyokkE/qT5uCS4eep/1jPQqC6tSUCzaqPTGUADgXD
VWYj1uNLHdO0cSitUsygcc7PcSqomQs8luDdkC8p1ua1fEA4EHNOAw9/o5pEbbKW
YLQlYaM2bNemvgU4Y9HWu9YxF+LvW3XeznmO/4CAOb9fr3b7vdtfMjMgAQHVmgXD
qOih475/zN7S6nCzCcTsjFcL4kOj6rX5fSxqcJkudU2K62iUDsekLn9NC1S/0Nm0
ycI0woY+K53kZll6IpvLhP8qQ1fmvX2qfDBxPZANOcp0E80sSPm1Z+257GtwIgfn
9SdqKj9HjSsj7OswL2DkUuMfv63CNDbrJ2z9Rwzs83r1zSvdmd6/4N3VG2x6RTeW
09oAQT+wu4eT6yKMz1Gj1PVdbpiUZKZ2lP7L6ca9eIyYZEYGrDJXOPc3C09Ymxc6
dON/0l3fGFiFSS2P1KzSzFmAXAXOr99jzICbw2QuFUPJesAYUuIp4F6odC5CNY8E
7Rgy0YUffprTmOuz58eIAfMxDUgopm87WAinMXn4lTawSrvJRJt2EJ+pkTp9WXIX
1FWu678poTTqh7D35AA861vKK/IgPaMnQuXoKUn0JeQ0v+aSQSCNA7rKir8JCSnu
Q61JIF3zqzqnrp34aiGxYbz504alOpOJVZPHktnYX71WUxP6K2LkGwhlGe5PGMqx
nk9ZdObR7746dZrBJFga2hZbeqpFj5dj7udLAvKXRxUDuT8+1sqpxy/HqVWH9whp
5oAGS9JsEys9L23pxKVyE4HcLEK8B/ssFQQOY1mqhJpniCUIbPXtLRNJMaIF4erE
UinKs8cJ/ioa2uR4RflOT44rmVMqTx8zaYzYNQPyA1PS0c855U30JOTMlw7F8S/Q
ZyaSrqgEuBc/qakY2WVbpNUdwAOBscr5AMZ7ilT9qZ3DuM0v+i8v44/4L2aH6a+s
bGjvjOuN/KuzE5JJ3hmoWMRJ7vIZq2GCV4KC8kaed7l9TpiLf+6PBG7DuooFx0RZ
p25gJtQUNmXzWzn8YhwNTGCYCib9sh2O8uMBi1KoqpIIPjDxlba+uDcLq5r60zG+
56C7Qnd+UD9r1CGnlNjzCPLXW+yYOLloi2mA1FrD2UoDNYNtTEZ5TPlWH0TxYAT0
vk5d3HynIsxhIYANDxEkSrG4xnItUnctUE2+cZschSt5ZfpAfOzYvowRFKA+dqa+
Iv4ZaATErwKtuQPPL89CfWBRvhymCq3CtJPc3erYwyiK4fXHQIZEGiaOL1PUJtSS
t8VpQCdzs6U7/MbBffK60wipWIuqIVhxmS3L3RkQ1a6kCuUu0Dxw/jzww8kPcMfg
/nDYq2QBYrFmukMopfiDnkHMoqNuUhHds7yYJSP3lwmHlWIsPNv3leFYbdt+BoOF
xtSVPRfkIP1XPKodWjB4/0pJEkBu2Bvo/1GEA7Ep/eV9lwY9Wn/xs/HseQyyCg7D
eV2so9A1SWn77P01UEhQeGlzo+YXFfIij3V/hu8jB3HIeVi9tV5aMFX73SYBq5vf
BRSePFrt6nT9OQN049P0AbrPx0n30miak/NJhJsaFn8Ko04P+aE9QYAbz8MeMSzX
7dQ212nLkZeR9UYsi0A6JNP7j/lXV/ZEm7WbePEXASq1YH3hps+u3Hj80hRZfMLp
mfad5Lply+ZM+yNrSdO1L12TxlW4VEWjl+ZrdHQCRG9WvqRacf5RjtnOa5VQCdNc
pvgW/SaryEmd8HoHevENP8mR76hDPECQut9sJs0zaJeQS+LdTzcYsC3167x70HAB
9h+o7Zu4IXVn6fVGanLMHuyXTAv/YGDdNx5w8Hf+Fv+Wxl39lppfQPl9stIisxKE
jtA/ou0rubcwfELeXeuLM7b3g0ZqSFiP8TJiSRPRFtMmgkmHxp7pn/sqEsVXjIrG
LCW8lT9xwdtOjo0yGMdFcLtQYJhRBqC26nc55jn46miq69sp3RH49G1pUjjh4kOJ
JMqSYXVAw8qk+ExK1uuD5O1DHuakdlX58b8olqXhNiASoXiK0TueMZQuMHtLJfj5
zcuhGbF/rVKIuxttDe+g2m7T+OCHqg9EjpvwvgdWauYlRp8+msjVvT1gs99FXf+N
Svci1roINRmsvg/vA97WKBP3x6yxM0EM2HgzXWs4tF+Zmmzyf0VPE802l42+7Xzq
1u+z12JeOhGAG9NOG5p9kLePPZ6Yj6iwKXzFDKX8Avxok7kdkGREM3ziPq328PRC
m23y6//bCvfWg+7UcwM0V4kZfSt0LBx6VzPLj/EbkeHpW0TkAXuU6z+BqJ7mTw4H
VMgvDSPfhBk/ezPagweGdfWrRoGneut9poQFmFouVkoko8/e3GXZ/muq8IdjeYHH
h5yhtwsQIPUt0qjh/+hWewUwDxA44Wrei+gJD8VzoesY0AwP7lO8Qbv2KFG389cM
fv51Y4WQb4RBrX/3sV3wMdT9qcZCmTP5GpEo/WK366H7mAIQjrLOffRKF5MU7lEY
cHM19+grPvZCi1LH0M12LD+KMJIklWG08Gkj9ABXMfAivVcqBMZIx95ZsnJVj81Z
UpDOmsxUFFTbh9Q+iDxxu5SHxy6ICL8/qDqPqbdlLSXgzJrTG8Bgx8WnrtGlSIiM
YOA49u33Cwbi0csbAWR1sDtlWQc4tB1GBZRfTMI4JD3IGY9pZICY1JPZ9gGE0iTi
43Cxn1CbsRIefK134UJp4oS4Jzqof25xFgkQEGa3yAbLCVufZiiBsvOemALys+je
NyADrg7tA+hOKfFiYLWi32hFUOzO68YDyh6d0gq+fryGE2gIPyITRlbDGNCSOrXY
B1wMqU2YSf780lJ/TIF+iBwWj5xbhAH1q1eyGrI+KqirdKy9sLBsHS6DfuF7k/qe
hQlhTar3FOwYZ8vYJKPHiwIRPfztHlxmkUgpcnTnUYeqd4wnfcnxseXNSkE1l2Aa
zEI7Fx8hiJumvzaP6un/1mcMqb5s2pWxyNHhzVeRZFxj1QCaw+nPtcWxxlKssZHI
3yZScWH7UIIOnUoUwp6ShLW2f+rrCYDgmBSRxzbZTbI+eQAK9qC2eoroiAH7eIEq
CiEqba8tQiTaguw3SZ7vyANI8utn99RBQuYwaJCwhIt7/lTr8C3dV96wSw5+0A2s
09YGcwuBj9ssddRPKV4AO8fSLyN6VN85/93yf5wjOdrx1+w3x74A7YxfRaEeWChX
fqGlp8jaGFHOYt1X9Sg3f8AAKHUzqIyHaqqmpwluMt7NH7JICyG9n0IJxkC+fj83
pHoX/qzKY3aaXKj9LF0dpKsMdxiJAShAGBODyw2GsQ08PmgsoLNqQ2HpMjjCsFhM
1qQnK0NL8fs3L4kApkLcj5G83woqpQZuhRfrKEstqkdHQiEUx/qgyRYy5WkncD0C
yqeiikMKVl7eZgtZ7CvBnZ2yELGYZCCTxlT0B1/GzxTevyi2cqNPKE6eV7d8k2Qp
QJGOs2rtGnZCM9vu60kam2zwcl0G0jypxIVMSBtMdsc1kbAcrztpWagYa1oozXG4
bA+q/VlDffcoH85SJxdpQJcOWXgWjI+jMoQZC/oEZSP6x28Pp2CnkMh/eKzaCQWC
SwKDHAFjJYG49Z8BKyOBn8IQpA/vovD7Oma3cwskH1Uf4A+lB5LCVs+prfDdJ+V5
N9AWWc8Fb/7swMt0Ct5iyygXK9i3875Qn061auwaYU8guSrlpExaDLHhwkRIQya3
JxHwUhAh42+6/kg5Jhc+Hfhx7Q/LAN17EpIYCQJs2DQnd6mKjMpzi2EcfSOsjXzP
VeyyNZx8mE2DzgbTKDAQhV1vSXsbFns7MXiBbLpcgBaoxq3EESf2qeyWJdV+6aIZ
N/QqUk8a1wGii+bC6wbEh0k3lAz1xEa8E1/cMMAiH/ANtOSrX/w9gsxX3i8/G7Dr
9gxZ77493SPqZfY/Yj2OFI4dH5Hd5st7M/xxJqxGR8ZBG17B/rZ7qbbl3G9nTe0t
MOd9CVIWheWRCK8e17Msu7Ctqf8iK2bKSe/Wp2vJpwGVEVgVio1+MEk2AC74I8co
z9yIml4c8lCkd6RPmHhGngtqTA0YoeIGfF9hfRqTZlglbWQXPDOdLKA7MbYqv1Cs
+99RtHBkGf1+MTBFTxzmA3zgwod7K6coc0ap79HUDoxDsLkcyMwUoUA9EV3RfQb+
r0iWAe748YrxdOVaUc10LdHkOWzd2brv6oMuliiAVjzJkHENMoM9ehwTQL+C8r/2
6VZJ8iAfTwSL55HbTMHnqy6hqHZJFgNf28cjg83TRTI4D6vDb+KMfplHmXEIwrA8
dMpvwmFVvzlwi3PxvqHZsrZtv2KR7r3/gYpAJ/yp70y+ieAOdnTcLoqZ4h2i7bhD
jOE0vaM7D2Q9kE4SnVAr1nbu1RLS/94U9w6yKm12xtppDvbrfmpCgLPF0hjzUuxG
LzHe1nUyQkr0XrXN5VHVa5MNiTSkvIm+q4fikMR1igzoDbHpyjLIMk5PDm1cp3UG
gYgOzkQu8aUsULr9G+qf7aWBjWM+f5GkxEYmLqfXXjchbbhWEb3rgyheBu3mNWFH
GMCpFXSaXhVi4zgXxplERQxuznDMN6iryGUu9GO67idDs+MkphtoGTLPEOs9o3k5
mwPaky/f+fvoSAsAlbzdY5R6BkZwRjjj1j0aQtgU4UCJ7iiWrd7t57cHo/POPCwV
et2PB8tQOiQbA77lFwMwKPzhO0HRBRhe5AqJUt7nISE4KTlt14xtD0iC1f9ErSlM
eXv7qyx5WQOLkg/GhDmg2VIgiUsQmtOjZkYp1oCYeAJS4NYQet+NqvReiyCcW90a
Dv5zy6MRLb00K2KP0fFDb74FqxFalIVcpimafKtZbtRx5vKFL5O2M68DFhF+C/LO
uJVqIOsROEmNrY7jbR9uTYjFqJLtwlxU93VLLYQ9PjelUhApMWwL5fB8vPXqwva1
qTe9aqNtSydH3bxyGaA6xqcFTUfgcbyg/P8X2x+3JnytEcspuwrOmWkW4jzbMYvB
fNbDtCgq54L4ohgqCOkkaNNsCW0deotevg8bPeHD/czmRsY3Q1Nn9buRmoJOD/jd
hy0wru/nt4s/GMqWUqY+J1iNBGOyXy9GrKNOeCg5x6TsyJPE2QbdA+y5ws4q1xPk
1Nbf5c3ASUvbJoTLzi5Y2yaJVhc5xml7NlXEs+N5cNJ8tVP50efPeigWvYfrbwdi
9J241qudWAfkbD0nEd153PeAK6TmyaPPX9BYaUKSziuwlZ24jWYYvITlSIEJhWP5
6qweJenD/o/xm8kZlupbhaditKlc9dQMAuS/mLreYxfygr+iJfy7pnZ4qZa5P1XA
9+hG0luskVgPlXn70e+CVdgu5Z4Fp8eClV6t2e3+G5d1M69h9ZRtS1FZ7Mmdcp6q
76Txq5BzICoMIj7ovg5zXci4wFfnaGPVWCUheEz7NqSf+uSp+Nt3TT0ExVO6H+lA
Wvi4bgGI/WrWFg3bWJY8eLYKeHfd6zVt0fLt8/P6uD+ggtmXMtkYedRmDyQ2diL9
zVlSrHLN0p1kJsUCO11oI/izIqSeryFOX4Asj77luBM0oN43SipVZXKEgx+dB/Om
is1+QcIT4FoPoiL52vu+QRfB+Af35odKdzvilTkGkI7dAMb40+diOCmKDYmLqHbE
htJXfxGx/wiM1LY5LpB5HADAF0f2WB03F8iwshjDqGwkLpXKKq4hvndkidqHPRrD
wDpoFv8NT7KMl1YuDM2D1i2tcrqEC88SdVro+bgauG9Xn/BxUbvQxuFbT38jjF3m
uAER9g0KvbAecaFZYfa2DRkP4SmdAtNeF5zA6xv5eV7IUHkLfwcdamx6pQRtFPZr
QPPiPxZeZUe7QFKNQI+RI3j/lnaJG3czeriRqtT/Y+OBe+TwyVvDJ8wCGc7uekqE
1itV/SN/GQDpxAmUvPebTbhFSwyzt+VTJGfwIoz76xa8JeKT39b17TRu27hBXSjA
k+CUZrOfPmU0ztHXzUATZtybwquySLcWW4Crt9MqYpgKxHA5u2E5+oyONhS7/543
4xKAikeCEEvm8IsRT1c7TKrOj+dFAtfZ37lnfdhz5Mvr2rFEAHpGrSw0KY+VnIJf
ZuiFjIWEl37ok7PyxQqPrxvGXnYAaBFMLoXjak+SCRz8VfqlRfYic62Glwf2/MDf
sG1Go91Kg15H43y+s+h1AD3UAMtKs8NOKxsVEpCf/KTd0F+vJW1cgGyeCjVjQ9KY
Y8LopfJfUB6dPOOxGncjcuVrlkAE2cAVMWdFm2AbM//npdGG+H67qlcxYpV6evU9
kgM7sPPEef3HjS0M8wLzbLfA/zPKZOXxy383wDMi5JAW94prpqWLLvqbdsm76eYi
dSiMvTy+KBh63iIo3tV01pq8ePSSUd+/SaZ9Zia07x2osbLU9O0qIaCsklkZZ4XI
QZyohgAVLugu1BljbZzLsLTMjEJiu8Nscg+9kNDy0gJoe/e98M48noKUFLdL/29A
E+EbTQHtkdE6RGXP3Lt5A4SuqPQ7WWuZ8eUdK2li5UdU14rSjn5W6Y2LE1by72Fz
lQDd0rDaMqnYhpGBuQLiZMpyCUcdiSIjEYd6QNZzW5IgVPKJ5vHwv2tF/iRXa7DC
u7JGj4W8E8FkuuFbYcAdHi4YdKSVHfSdVwQE6tn7aDaNdJ+LoU6HTuDum3NL1T9H
ptGkC5jW1gcyvS2hb9oBUhQusQtIFrES7qTIne492j6euY9zgn5vHHqQj5kZfeXk
TKWZkk7fQlNeweCpmw3+ysaZPLutr37SGARLPckU868fnOB2VuH6CMQqwPEjWJZ2
ru32fv0pS9k7KXhouhhuqrgEeY6C+3O063Iv4Tk6h6QsQKEGkkU9xVUZ0/JGwqN+
LOZrt4XcFUTiUdwlViLZQoBGMeetiJCMhw9fPa1RIsuzka2hSd3WQI2OZy+ofG4n
b9MAcCfUW2g5UjoY+ANd3hiVg4mipDtoZ2c+Htdrs/Igw9KNgk8kjGC0u8lcfzu6
++CYOgR+I9ajmQRRpVv1oYU51BaGzc/fuRP84vgy/OVDoGCJL2lijFbpFfMM48fr
XBjU3aGRLXsehaRs018GkqXwBCmF8bZSMIJq30Dy04UEqJ6esWc+YA3Vf4sQmXPx
NVLgWUF0gb7R/48WV3DqXAihnRXoqvIzj8f166Jfj0w6a3VKUTYkpvRNaHuIz5Jb
ufOXWOP6vVzNjiv5UIYw/pzrqjHjxliCdvwzBtf8rwVJWlNKBUWsl4qvORjQqXQ+
B4H+Y/6p8J452mXaATTyuYYfBuA60K1XFpf2cQO6OYlcT1MtAOxPR5y2mIacMv7F
LmTFrRVPNe/1MilEnY0PuNFqQg61ymqtgIKoa/uwxCOyts0COuB+Jt8PKk/U8DWs
K0kq+Qh+Rqwu0pFHqZa3DVQgyN/trI74qREjBnDf0mEDRqeHJFxvGFxo06OQaLRr
09nD3sKj1pTpAvBM8YrDmafJAn49/yYs0S6u7Vo6a0Cw0KSQiMOzPVPGnBTHomDy
fhu0KgA/0/zQZxxEZYCD3wZA1DhH3uV6mcEgkGcztFzJgFVMVy3ZtDRdrb9bcCAt
EyUtvZyaSVpebQqlX80o1LnfzOmzSFM7vdVF3ejOVXXphIP87KxQppriJAM7uS6h
uf4ucgiC+0fkDaStx798HFLajx0daF9coHurIwKjUMlmOP808DtHVsLK1VTO2Klk
jIyaC+3KYL+QrT038/W3kSfJHH6/eYMvynqE+giRf14XCSoA5lp1y69HEUQy6lyk
RaYjaKIb9IRh+Oy7fC3OIMzkvmKW6cPf1v3VYRco4N5oVe2V6HwUqEXspteQT6OV
9rGzUkMHoq2wxbr34+YXfv1X7h7RBpk1BFXkjX+t4AU+zvQsR6v+Rgjul3wUsFQ3
po9DXHO2AG2npCAtmoJxyMObxRQzCPLQ6lbojIlNsohRqF2kNW+rJGTNLMMOIjGg
OP9elZjCeNzSLSWVo7OfsrMCcosw1+uyE0HrdqB9Rer94LFpRo75ljZy8GlXh62n
1yWJuTcZoiJE0vw0ZuPlBeNg8rFAuihBqP26BxQqlNQErNRbswwYuyHCytD1B8V6
j/UppYYTk2LBtWoduVc3CwtaZmlvIXdz793qpMETYnQdAUlvtHluvnQ5gTFy9CPz
znzSaHxRrp58I1Tl3nTUcDF63llC6jkUgrY1+tTdkJI00i6F3Sa3SHDcwilKFF0h
UahiZkqNki9w4Awt77woroppCJZQHcPO/+s+iIJ836mRfkta3Op/zYk1ssJymhCy
PC64e3Hwls+nrqR6BMvh8R0YQ9WIReu5recCtbgsS7QrRyhJzHZ+8pDxG/NWOHdv
ePiUVmZh7v8tg7oWISZl724eTqbD4dTDvpoluGWgDicRmVavbdQcn28oAed18qy2
xMEG6YbzDts/gbRC03Vk0jvdioFYTZgd5R5MylUbNnCiVTJvjkLuqVhhDkUiA33n
1HuLwy0PIwy8LUKP8dkBaookkdmBE7Xb7hDazo+i+VVkdLtu9OPZ3pIQiJOpFeq8
TZlvAgwtuoczpJPxWXJ00oYWcorkOPTF3bOQNFro0WcQPwaTllWRdgj8CJjBavB7
KFrd9VLxUZkIwz33NDQhXAwNL9Pr9UULyIO0Z8R55ETvzg9rdaPU5BZmc+/c6vtY
/sVG1ICCOrEUvz480oMpZbeR7MOhq2epS4B9XovpZ7ThkrELgFpGIyCNjCfjUwXy
0GOT96Me7CpXDtAntIT+iDmc1F3atcAaavjtH7ARVCBKNNQUSB3ZRYRIXzASqyDc
/Zsspr8axXiB0qjjKoVn+H3VY1l1Vwn10JomvvA64HLa8KNECzwpv8pO9P1atqKM
duFUuQc7lAx/pV0PsJKrT07RONwAlQke/ifunW8AzzUMUZTLij/Go1f8JjHMGdZk
L9fmoQSXvLTgFSQeFHC7luwuzpTGxfmru0X8s9TuRZI7Lnwk0cH4mKhBRAO3fBr5
5ic4l16Zx3mkr9ZbKNX8yo+aSWfyAdaecF22GG5/6yce+0OBTfxfSYdvZISzbJXe
qV+goJjr/HvuYZJtfZsVFZyj436VTTtD0lpix5L2Ef/xHNyLXE9teBZhSutI6fPE
q2Oz747dib/SnMfRr+cQVRotyIy+JTYDNcqKGHDseHhm5uun9dBGjUdzPbNP/D5A
Xrq5oh3LnPJMm3kVEFIKcMc4yjI/tUcHAqmOdwKPjXMpuYbkm9eTOniKIZlBv9gD
14BoCxHIjiCK3RiWnWy1SkqApharx7cgsbCixw/mfYh/rNTqZh2QKInYNmrftSkX
0zyJV1y8sXls0UGi9CjyN76RKjSrCulSuyq7rV3uFZKCCVC4dWzTsqzn7ENtaIso
9s/8FwV/if06iAzN+KOiMXVSGdI54ti2IeRjmC41maEnQk8T05hpWQhhsvyQmOcv
z/CWfL7Nh+zfmbK2eLOXi0WUqln53U0nVjno8hZD8QrvmmnokiwuRGa6vn3DkJES
+g3Npl+KhzC9enJub73ZybYd3vfKCUgUJnwhuRcckO44hzA5DSY/6efnK0Vf8ndG
1/UMlShOWy7L8pjiuE8UdmbKVC3QUAjq4lHjEsc7ReY2rvC82H1aRPh8QRuTs+ff
8eBfMxmQ77+luBe/pzfKXxdnSgKFpJyomK3qi1tNPb3WUifAA4RFNztk1haG603j
PRCGEXrdlaeXSf8Lpct1UOnbvIbjoQV0RapUi0uBRs3eMLgvlCh5CRIvx6zZ9XfT
LtH3ZuLiKazmL1QPHZ/sfGaHsog7rD2vS99anwjTeio3ICPhQTFZGHVTi1jYhXFs
OX13zlOVTIXpPbtjuFqR4uzLgkpSDC1Q3H0+yn3A74FFzgdtOboMU7OFHZzJxp4m
Ajg9ocefIem3e9D8YYKK8fARsyKsTwqZS0F+1JL7hZtftfiFd/exejm6299GqYjn
j3x7xE5nzuGv2LJKJZb5Xy8SBzgX8q0uXsbbixFD//lnlBDt7Bbs/iQ3AjJpw1jo
6fszQmdEmmI3+jNhNOfG1DuIc4mTMPditOzEHMkdqHNmrf3aoXqWu17Qn5kTBbDu
EAd+NVLk/LtJcfaiG6n8UT6Nyx5pX4zehtJzotwR9uIVXfEe0A87Uyseab4Q8RJN
DakiYZBqvzrhIeantd4w/dQOOwFy+AMaQRudJ9mmQFDjxEtK592Vevhd7pUy8t0l
UlpsOSjM2pCNHzAsfKPJwvhTvRA5hilThf/B+12cTJYPB3RH1NUZ+1Ssm/jQh8ZB
BoM26b+qPOxK6wMSWVTne9kGGIh7C29I9cxaihY8m1ZTIUK8CLefDHa4WbTO/9vm
PmwohwdlwMX6GaH9O2/WQOKqmjesjKM3aAMS2HnTCD5dXr1KvuMQvD8EALqK0N3G
Lx2z4MC3+rPcZJ/VbD1+xIZfhnDr88w72wQgUWYdueL3Y2p5e5BJs4Nmn2y+4D5Z
BPg1szK9vD5pSlhmsbeaqQSZ6D12WKszogjBqjgl/stOi700LotxvJJzQBfmkxLC
v7nTNHrQg/pl0M6aYmKtL8ONIk9n06N1HKotsAMBsGcIABS5SyNcCKpubIFC36DI
ZoB+NmAZBpYVJtTyRVS4N5TaLICQjBOAhjSNEIFq81dzHqbVKyDtzgu5N7FXd+ZM
f5bfongzQza6a1bpDyS4ybtbrpptKQAnrKeyozgTsct7Dp8f/JpOA80MqwI87Iup
F6ee7xKwjw3wriI+w6LOhZkBAfSkDX5C/Pz7lSMaKUqsyBLULofM+0awWNASq2rg
6HdK4B97Q45Il9Fly6uYxv+Ch1KMfESQQwn/URAk3HQ+sDRzPT9MgI52yM2S+GyV
FU7jUrtJJTnoDeJs1T2bd4FkBiQ0t9zD0u3Op6yuzMYRRepbgEMEW4w2a36X1hDk
UIyqSqIY3UTyTBUiRZsGQ1zPlgyAB2lCVQuei32kNlfaoMFFJINkvQL7WFdUUq4o
NsBxKy3WA9AuNGqDkXMe4RcE7FiCCSb36hEO7fpeMqP5zrjqAK1J0X3bG8XMOxPV
ndSghxBUWrzBvbgMguy4UbEKY4Ff8Z1MM8EArXYB2OTZM6F46cvnuz0E755SaPoU
0+Sj+4lRwUc/x0teEo30vP0ApjhAE7SPQO3yEXIQjOZdw7ik1ZD+V06W8/nPC8Fe
Twt++GsPAXWCbc+2GEjeELwbEAhCJWZwft7ZxIjIsbO0KlT3CUUQzyKrECR5ifFB
okrVhM7REMToLJGF8q4ymAUMYiHdy8otOKngICmznbEcUL1SzCxSrD5oLqJ1iVUJ
7KlaFwe0InneB+ydAT2jo4A5gyvkmV4UAHdJRorlLd2sMG3EDRNcchrNLKXuJdBN
VQYKkN/J3f55rqOk6p28NnpWISdj8EwX9Lx2CXh3LJihxWO5Lo9xJrm2QnKyAZX6
uNAlEGPtEyAkUOt91/C4otXov3ogDwwthhlvYrNusIHjNroRgNHvCJWFJEdF8dRQ
S3qG0I5RxTxR/lQ0dD4ENZ4e1maDp3NA5kmp4knsEZk7+0VoY8GnWZVDQcbm/l3F
WuqdZD5IOOTPL6wYVgOzJI9K5fEaQpRWGot2sLa96yLIsU825LvZl8mrHEK38jkZ
HHS7sT3s0JatyGN3ElcvgtG08+1yvg5Mt3+i5EZ/tp6qlADSaVSTnPH7t9RqeKEr
zZHNnmLE2mwC3f3JXIgFpA+h0Vt39+/VhmUUz1JFeBSNfxiWfmFfTnpyJqQ/nrF8
VEgqyTJsJsWW9KXEumkem34nmbTudgDkM8eRM/aUTg+0G0oCWMlYYTN0ZdVaVCHc
KUb7lcTYTbZ0FDOhvJElJDzZrboL101aX8kw2T2mJdQN2vApYEPiC1o0oUA2B7Qa
3ctFnx1Lj1PJzleTZISdztlXg51AOOK11TljrohUhTiOXaVCcpJJ8vX/AU34P+Gv
yWaQezMw9NnrQ6ybGY+G62smsBKdfQCNdjIaM7HO9H491lQVvjuKK2kFJFBKdof7
K/a3jfvR2KvdKRDZYkW+NKxQqvzDx12882sIwrgr1F+nVdO/YtF+PhA+mTJ1Vsum
A1V/htqEP4NBdWH/VXtPJlEtaMBj+w99n3Mq/w6kh364qtNmwlFekG5oxL6/eTqS
pZYteApodZ5QvcOEMlqnm5MCc9kbpu8gAcdTCyqB/SawmAYjKAsxVZPB4nPJLiiC
z/7VtYnetRqZ0npRhHFW1lyN6E06FltCSI3MLvnPeOVOhiB+E0w5OOKAA0GDJPgZ
LUn37mQEprQ8PGc3v+R+BpQybWMHN4BSZGVNeCv5NqLfuRf/DlwHvGC7cko7Sfbp
UIaMkL638IyRyo9nnIMq+r+3SqdBq/IbVV/HVWZtHu/hFPGHlTW1IVFOfEwCBNmT
hbrPOh3eLanFKxdxrKDVXhRKGrm/buNvjOAP55GFh06SzDAApuF2vRoeMdzfxpKA
0Ev5C8oM4Et/w8lvKuXtiFNMISoTfRUER58UE5B7pXfJDr5p2iY/pIIXRw67jWga
yYGvtZJ/SOMMlwbDY5CA1bUv7SbvSI7QA4w298IbHaw6/fJUGU5N/U8/lzsl1O00
F1+2FdzIH4/Bx795FTxTxR96KM9M1KddOsl7Y7UzbLIXHrU5Imy0b8CWQFWP705G
uSLt2ItZefDrKTmGcZUa7TrK3BmYdLlGXKPnvLRCeuSxDJfUrYUtQJoHkBoeNeru
3moZfiovmvBRLLQOEU0lYaSqz6ifFWTMXvbDBzjNSXYuTnud4h67xasFXD0t61wq
Xbg87sjL9EBEN9FiXerUtZhEJBIbap/uqOu+BgUBEhdavnBwR+QXHucMbSfHUfqy
lOdRzCM5L+SGdMhSsVrSD2R/VaJOjFwHwNinmr4+Uy69agUhVVqf9967ngExEyIv
PSUCQo3UqXgRnD05/cUx9Be7jOieS487JxLJYefB/YxOZuORJPwmM9Vj2tq1vcdO
+oWGWhKQeRDwmDBehmCuSC1y+J9pN4zg5QYHDy6/CqONrwTu6jIBJYJpfFIi73Np
yr9urWwrM/lChqlCU1n64vs2PhT/MnRDMzYhFk/YsqtmakKAwshIXAKxiASZy8/B
agNkSiNdybQvYsw8hpfyjn3xVBaaLuDKABFRgaml2J00yeU3y7cDhWNGPE9n2u0a
xApKVpA6XJevk0GsM0/5PtxYa2oveg1zf9TcczjPsKM8lmLJaJ8YRjIL7IbCUzWT
GjFVL2XxDROd5SQ97s9KBDM2cgV623Ax2RlLmCUk80KNybPyLtcnLaNT3041QHQE
flTmyVOBFPPnu1KPWBwaQe2xcWwdk57GRdPKscR2yvuvoM8Zvx/TM09uzpUJtmMe
t6/K04NUMWoEPtZd5N4InKALX92qrxlFv/wKmsr/EB9SEKdxQNT4wEfwum/bnS6k
uXKxIIzLaClybAHo4kTL3FsbuXDLsB0SW4dYYQPN/A7tZy/zkqQboZwvJMMxnYa2
Mpq57Wr7IgNkGDwuQEjykPElNZ5bwkDzHIivAK+NoyBn6qxPdmzPCAj5B8sUVX2c
PX0MoCZp9lFHkq0ilutWitgjqEu3bz3LkCoZfHdcVuJhQlFbmA6da8/qiU+5YNaQ
QrngQE2fQw8UvEe3iUTebJ2B2AgXN8d2IphP1032qSqZZrquKNyWDIL9XqmV23Rb
R7+/wYvg1EbKHJpm3g4kqZXswPM+uRrd0Ugu3zvytG7oCkfdsyFv4x/37CfxFrlN
kC943E93E2O1eMzWkExE8kBoq5u8GaWwLFrzio82A5HIKcrL0hwKGrxjhqeDAPNe
iWOEJ9XpAWUDLySYAKeUuZ2OEwiJpTkCzxjxHpnFn50AKfpIv5QGmruN+iz463IE
HF+CkzJPJD9M1IHhDAwsFtqWtTbeeExXO7/mOo55+/eXqT2SQFajh+X5kzMOjQNP
qpjRIQQ41aZW68mF0jAPlbufIlKQI4QPWLJP1cvXoULcdMzNNtvjDhT5f8rgA8XX
ru57B/MJ+z3hSwu8yagn/Al9WKzpFBbxDsH/L4tTyMTVVqeOuPXyIpP8VkgofJNO
E4cCi1a7v0fwLX/F3dYamOnDBxbAlNauMGEL475k7YdczzZ/2opmyLpwn3l0eBUl
ejZK3vNQkWgzmro1p/e3fZ1mJBOWpMQ0uZrRiAePOQaitC5Fwp8EV7B7fplX8Iwe
7XirUwNcjqLsRERRNIOUJRekE/6t3umUSCJdoOnTPZrLgrKJzpSWDcaPxBE+vFdp
u9ZjS1jz25mQHdZVhSA7saJsOJ5j2/oChpDbg+ypXkh/VZE2A5ft8FtSAtaLfSV+
1KC6sza+uzJRg0zbKYASI5816w+3OXpWYfCwuLUCkkDMLAYfDL56/RPzFa+VA3WB
6dbSi1iGrWsZ18DCVz8JF+8xCJ8rrrdq/SR1ldVUa5afw7qIk/u2XtfPZnfegs4I
kfTNksevmSEF8gSS4IlsRiU36SaGE/9IjkaMjjXpNYoasBDh0G2tP+E4Jn+oArOC
BlVebT3oty957T3zqbcOlEqYZBwol/B36Xz+BHu5hQcOCG0gkoMn46RljeQcw/7F
Tnlub4ViEOWuVmjlgQ5WhD+1zrqrZKMyRoO+UTpifZgpxiI9mpXQnPD+uA5//p+1
UN0DzYFWuJveLXNbsNEIa1pVf2BinL4aCCw+nZ31Wplhza1++DGWR4x/LrLm+W6J
xPfT/amWMHNyfMWP7CkJPmZzylLDdw2GPJZ+6kA11bbxOKhPtgMBwoob1WCdCA/i
KZ0+SJ7W4jvF6rY3sfGBQ6ANZ9OUiA9qNGjFQ/ygIv0gd+nWMkCADG2OqLGvDZrp
5X0Knq9Sfl3adlpfjIQFtfWwh7DvHhS23rtu3Z/h9iG4X+qhLCzuuQjPNJ89kpFx
ul96n8npxw7KQhb85yzPoAD12uuAElQhNB6b5EZ2rdRFdOwoFotqN9yABKQbFur7
srCbgdu24edK3jao3kL32uRxPXP7jtjy3Q67DY5yFy6/C9EnOryln6oJ/Bqw9d80
gxuVs/cFk5XbYfBCmCgh6h3Nd/STvb74zRjWkV/fJTiu/KgJg6EmYevG/OBqJFsf
J7xWDIJ2cZaObjV6RZF6Zj2cniIcwLuEsjd+EMHauZX6juvxJgni+mkj/hR7yqJL
HGbPvyaRltdTYIf7zmcQMVZFZaOAuattnfusO88T0S7d/4wwXO9e3M5DoNliQAEF
xHCPwuF9fzhn0tLbNgJwSpyaUjvHLzXD/mEnF8tmlS3kayJKF/OGCoArpPhKwGVs
HkwbzL/dL0BYEylTaPhXuvxP2ekR1QBTJnQ8xO0jLdvbeGqeQIuDSaJtJrejIDKx
r/9LXnl2paVn5W17B1fBP4EqhExBgC2UHWnEHGPzYqBftkWOoDcchwmDj9qfp2/Z
rRocRlWhDyepxVPG2MBu6YRhL7XnIR29VgHU5ho3yLBxkosG4QIbaktDGDWqpigw
CA9CKKpyV49NPadHDdFm77K620FDImrv0ZNiN9/5lmgTQVOvfoowIcuJ0SRCq4Zd
w615tQK7WU5f+PFqeD2fiPVHTJsKF0L7JHsl6l6W0bP9PxYAKlKpy7WrAzWtymJb
MQWadFSi6GVgp/FDnygPP+TqUBO3gZWXzqwbkQ7HhqRN7fXFGK6ft3w/0up6bxMd
vusxp5/PA3A4OrhvznIVsdWdL5toTASMjW9xYd6il7QM/5sg3Jb92ypq7x2G6GDO
aT/WZGjqqk4DG/CXoW9Nq1Afq3nRKFvuxBaKsf35Ew/EOIXXWP97tG7riLYBM4SD
0Z7Z8PE59zbNodym1MWiy/OD7injitBylRu/F3wZms+aIkPFSNSt/YoADAODyK+6
YzaSeNicT2XYz9yIRmLFbBIxlFUozLKHFOU+yoUsAs0GLkhUK3clisj56eY1cuyL
w0pP1Y432oyCfSNqmm3rRvAxoo68qvsz0M1CfMTGdda/s64bNWvFsAlZa09VNcBm
YIIxNdQvdyDdEXHsVubkZ3u21fCeTHRG2vyUGDoEwJXvqVH9twvnzfkKP19bHb+M
FiNGoEdHi045wQ/S+Q1rGKCI5ycKOeXquEo2JAQKcqNMPkW6qhaOKRDxLVs0suoF
8C72OMh3XKL9lkndySS1Qg1W77HUuTdSE86FPHPA+kQ/TgQ0PiDOJfUz4fd/WnW3
XowYEIqA7sAho8wqe9m05ALpdF7uqEcfswuH1WB/w9fIHzWxk+E6FO0qh4bppE35
gCK6x19pgk8qDIvHsunbIS8EDEdCcltmeRrLvMaVEof4fDntxsRteSfHrLKQlSLD
BzJiBuouEetVMOQW4dc0DJ0z0G1r7loh7Wm9d+ac82GEq4HBjv1LxfWLwxYcwwjW
ba2INC6cZWBHm/clTM3pdnIva22Goq8pVxGNgJ6nyY0/Q4Hv6PZSNf788t4lAJg5
DzoS5wQBoHtb0dbRaWF+Bii2F597DKucQBHeKTCoUOxpJwwoe7aDtcj+hlaE54Ac
jOz5k2pRFd9+fOR8L/OeCaGgDN8G3AZKhbUPtTclyJvnLF54jGtt2GvDLBzfyFs6
SWzZ/EDsIwkTvI7cWpzzq1h0YnZTgVHT/CKnbZlUfWZUbgsW3jmrS1VmpCJy+mcc
A9EZhkIfgh0u4LfacsK8geMtqssS7C6S+4af6+Mr4eAC7BQ+YCkj8zC3tCSIhvbW
j8AW1TJaOaXfHmjQnL6tciTaK+f31oqE6Bx3iizVi80HPVYzIGtwH9n/kydgh5vK
mRfyGL0xZnpKv4xoDbAXwabhHLzdM/Tndlht2l+RuA6xvOEzM9343mb2gtbq0BHg
QQ97JPBCBwXYwxRo6wkZFBNV9hEkpo1zWhLXvAn2iYhQEzg4y9OMDhjbcixme7ow
ngPUpWT5+NEYo4d8vAUNjTFQPPQbTiOl3XU6R2RfXHhP+OzpvfkTDYu4ghBxycNT
oUaaaFfTQ7LbR63o4yGUoRKQe+C197oxdXstnLu2XLc89xglcSR8EE4/Sh0AzaXC
gyPdK77Rhk/QwbdQ/pvuQa8xDMe1Kk2pR/OwyFPUy6NpiXU6NghM2a9gS3wOluO6
DHl9tkncfgZgr+VYjo1YFOSruQe31wMdr91KUleqM2LD2vBvud3AcXGxWH1y6hci
Z8hR19hJESxPkNS/von//vH3+vnLvBhkNRO2xr5IJp3FVM+burwlmQ9v+AawLTfm
iX3DcO53Xo/CKdby3jCUOyWkXD4n9s8+uQE0NvSE+kmqNn045PjsAODuXoZJ3b9o
VDJ9K4CgALoL67/Mk6cvpwNOw/ZRqN8eVWsYpUJSX+i/Te8udKDjZWJ6yDXxd0O+
Sb6tX7uUq+Lg9MDwyUgmhAKu5KPwmNGv39sEphr+UpmnP17fsFPqbIg/VwVxegtb
o6AAIKuEqffuUtSKanj7KpNxd4yU1EmZkrq0isrHxgZwjX3zsVP9mWQjAuvWQ9ts
rNXkJKt8gZe++VRtw0i1iD0O/fwHf+5o+GvL8a0phV5cNSQ0wG9BUY/+WAyUGwt/
iRMgOVJyYNFfdfcRZlw8rR/hE+D4KIwSahKMNhSRwIzGZmKh5UptXQP+8FDFlQgx
m3e8Plz19+9b8DRXcPX2vjHEW3KUCONF3XLV9cZuASkYY6jw2D0FTar9qeitseN1
Fwkz5d1sZVYHdUph1k2uEDLZpXNf4wAZBQcqJDNp9/uVYKYvnTdw87LHNnLCt5sK
bUbzhPy8xTNzmt5ksHRYS8q5PvaPJ3Q8KGrd+evGNfEvFOfz4oZohlk1/cjPLQ6e
INQRRe+3pUlNQ78pcLwzbYxQHk5+W9wohuvR9eUqkqFuxMhwNRnz49coXi9dChGR
u1+aWTkn8TP1hXHNr7YHqRxhzCwAnihRs8FI2EduyTf/WGZ4otidreKcVmetKR7V
J2L0WJBUkzEtRnLPgqutiMBeysj0E76ODKKboBBg8UDjxPUoAqKOEGVjrf3QGxRT
EZK0ZSh15505qRaVJ64nUZGLi42J0tRhkcFvvk4TTstmZgqwiR0WBWXFH+IA7BdO
gDzrexntoiU1yAvbGwT9ZZDmJzxyymNHBHxQMZ8KIHl7mTQcRe463X9mF8+RIx/g
t7cSZv2jm75eGa0VXhNAT5iRsJTDM664IX9744nBTDSR2APqulRIAmeyHmN3GLK4
TXRDTAWa7+txU5HllijrNxeOcT0AF5Gt9Z02qhmeIWb+p1cWnywssAaH8mZ/6WPn
LHmGZ7iitgr4srXvfOgLqufsoCthyUoDcs31tv06VOz22BfbFkpl8tnXy+ytVufx
SdyNVJ3MAeg+y2Q5P1VhFeOjfmHCqVEjzi3g5nTnSKyWawWbfcZDnuQqljYjyMGI
uQM/cRxV9HXGev6I7Xxho7XpTw2iQ8y/pI37KTzJ/Pzr7ThRiXkGDGfimvAETXLE
bTELcLgEQt1aPLU0AiB0+BPhTrk5CawqF5mltOcfoOCcZs9ZwrZNq8URXOw2pYEa
Wgwr8KQcdPNOAtDoeUMgpyXzIpBJZcZpl+0WIW35Hfx5Tl3QJjMjWGLrTQ5ugSw9
cgl/EMIVjb+EUibhZVoiZSS19niIUNdWcGTno2V2XVzrDfwb9+d999aTybjerqo6
i1t6Y9qK/IHLR0FhHpwsEaDWMHdoZI7D9NMOcupNmIPrhP+HSWJaQKm48mlfwsdg
CHMB7j67aydhhGnwxsfJeHAKNAAoblOYBMScwYTZUA/MBA03TKQxhcLn4uSLaKX5
gwN55nHRFmnvFLwgJgPErhl36NHUaiaXFKnSWxCrQmXL5FrpcOIz4tr9FetFdbvr
FFZQJAMWDKBRHMIEJ+eMUHszha9biXLVGi+XjSl2cfbFOHjtZeRHRHNclctAjUSA
tajzgXoZ3qS97VP6vROmtE7HNAA+PIJa0a6uTb39/pAyc6U1R8TkW10TeUNsCd0V
qxgzieXDpl0rFMQfmiDz0THweOGLDNXHmfF+APBe2W8JicfKMLRGVYED9vQIa8Gh
yDep5SM0z4wMbr/3hmYKUATcx+QAE3UCWVioNhmWBVSYZIqtbPQaoooWTZgNSFqv
NKkpBlaaCV+4PZzA69SzB6OeWTd+JdQjZVCZEdHg3VxdvuwlZfW4lvkZBGBeed7s
TLuvRKs9G4ZYTGkj6NqrhU3OETj5LTM3uiEGa8qhp0MB9PzJObE64mNUqJJl9a1b
tovDNvmBprgvtbhRppkZiZ27ZZcRh/9Nq3e60QyCuG9JzsQ0tmdrAhr1HSMwo5RY
uMLBB5Km73UzahImpa+M66H9GkxdIMzeVPvuURjaZXazBoSvKho5a3N7fT5n9vFH
hvRri/D6hT1tWHXyEKtS19ek9xES0qGz7rGsm2Z7nSzMAdK+WfyPZrJmCdNQU/fp
SRKBErgaidPWiZ8YOoooe3bRzRI3m5oVHTv/4bBB6NlgMIuLSRbfN7a0gSAwrdMB
yjaUtd6ARMjUyXOkLPqBtG+oHWV9KMNWHfEqN/0YXdGFbDKV25zjdh+e4bygxees
J8SHCVE5lJpAVJixT3pw7vwW9l6tpWGNFpsCOwPq7nuAKtErW+jtT3sViyuf/mcp
fMCUFLLTRN2k8W0/rj1/l92sIEX1vMo2nzGzsPVAzMWZLoxeZoYM1oFyMum9ePUC
d2iz4F5nktrYMUWmRG0Yr4THe5AlUo571dUHaGCSKc6TVQyof471at55SmiVNoKO
B1CEsH3yhBX+uosIrjQzL1mc8KNywHmo801yJjJGteJYX4wVH36fJ0qc1UjMO6/8
eX0D9KMXQSluLy+M/TblogiuL2NJOgBOVpX5zY1qcsYOiFuFPABvA4Y7CCv6WgRa
UnJ5t8sHdeky7OEYwh+ME2elkLBDdXHFenmfuYGZgXvfZJoHzZ3Sz86OQSjydYEW
FZEuF3p7ogS7l6ehRzOm3qOkeNZeduSbUiXE9zOJyKO0Ku7gm9aq1C1DWAha1yzQ
xNSLdNceD4lDSPkxxLb3GxBEUaCZwi5ZhUG+9Mto8UfDusPCiFw/qoDAkD6kze1S
GlX8h09U2FcMmZQd3vqQp6irB7jqu4ef0GMwTDtYAtMxsoGVHgXOv4UJE4zwheWJ
fJRQtuWYDnOluA3/usljXndBgBO+BPbvKflw5BeEdsqt+O/kDTXmfkr1loxoPo0t
3kTT6Q3wfvfNfvKDmqAQ74GHq9YYRvgNwB2GU/sRBWeTiTMxRWxm8HF1KMipowFl
HGZM6+cQx+OBxQqZJYg/0gNK4A25JOVlEPB4d2Yr2GlSRrpVi/5KSvpD0kvI6S06
eijDktQ4SP53WAb1fDgDcTHDjTtnFA/OQ4FoZVDtQ+DC2Cl3Gfr3XfETk/d8wFXC
QranYFJPgLTOxiLJdKIC5DubFmwk4/psRtzX1/mlufYTvtIUbgMGbyWRNKqLgg7a
pbF+QZU4HRlx/LbqKKHhq62lE+Qdz32aXpEyvaTt17tMhGO9QgJTlzLokOMDUcny
RKovn/ed6lgfpK/Tdzbj83kVksaEqxpQhVoURJFlTCTC3SuAYE04oavOloGSz/B8
XMDY18Irsvt4z+PCkbP1ylF9uRYnF1otYAzac5aXqjc2+5v2GqSlGxDiUuBxh2ez
FhBnkCnrTHLuV52ldlN0fQo1JAVXHASUsFHms6vZ74q9MmYZ42ge/Rfzgp+DBsPY
Ud8CfgOCdjOxEERwiVyJzgAuiMzERs4cWA/wCrfjT9Lz3GkUVEvg1um7XMmxcSHj
AbWQYP0L806NHVwJ33fgmcrNpDyAqfsCmpzTUYdYP7obfLWXEiCKLXY47RctBuzr
VQIxuGXPvR4IDX+h3jijavQJ64lbPXXO3X8CLq3nybBg/IFyWSRrH+MGzmnuGIlB
R/l/Y10x8bj+1MrsQcwwnUnt1pPCqEmqzkOYBMSwWytZbYlNC1uM/A8HfxqOmNUq
rRJnI3XRbh9y9N0eYA7KKWJjL6cy54U5UtlJgk8YzwXbYAnHHh406jpATZPwjSAY
e94oDrlibCgT3xc3ge/0/KaBNxMGSnkz2kDPPHLNG5xzJMi7leV7ZsbYm7nS5EKI
w4N2ZtKzfJEfUSbKJqesyudJXEMNAXZsrpmWSliEyBkk7IcofsaTjb4Nc3Mr0WIy
54bGOfQ/gP2tbyKGBCz7II/Udv+0/aeoB4S1v3tY3fHsM1xkHH72o+MVe+BcU2zh
bKoBpSrfLBIiSHQkGpM0qTvS437O2V6ipzVEFIHMpaKERcY7pQFQI25sQfV8yfcX
hlc+M7zXRA5TqL5+iTA1nrP0EhRY1tfZvkBW9ncMug3CiFMeNvehkksyN3Z6RSin
axP6e/m8JTg7+NQaTtZVigPK9OmPBO/jgLdXPIsNgG3FG5FIp3zXd2H1SmQjoNc5
A3PjQGmyZeq9a5KJqWx6cUW2pujttvc5wXXW7ysVt4Un1u7VwxNQzRAfBgBoBzIZ
ndRnhojl8YC5lAh+ZHNd+spQPV81gwI8WkgKrWDUZk6BtPwKRbqkT7v7CtlWeSGE
vcQn6FyNJnMt9t9kryH6MSluGoivl1oltL1RtlBXjPgqreAQrAme1VNFIJr+Ruq7
VSQggZN1gr3DEZNbgf5/aRtMZh88JFgQTzVvJkVUzLNJ/Zbsr8G2TaOF62DeD6yY
KeLae5CenSMzK9siCZBwS828tl/8YbbGPy8AMyz2aVNf0Q++UduOPWDFIxnjfK52
g9vfceOsXwuUKYP5IZ1hJbv5NF/2rdC/bK8zyfIKRK/S3AiQRdeKt56WZj8Arfev
p/336eeGQBCckkNlUbtEgiNVtInfjoeiju4XDFaaAeI/Pr5c6IvFWJep6UnEGDQr
/7nZhkrUJBCB1BodUQG9x+9q5gi7/YSnnuVz1mNMbYrDhDCrkqhmtC74gi3a8eCy
69MObuMv8DzEioYUfauAeOfFA0BPsf2+xgjhGwrKCeqv5BFtUCDQvRPYKrVwGfgj
RSateucIYbrsLgNWNMFtBXDrIDBNIA60le/KLYSrEnKmot1FsrYoTpon5ipPm+EJ
sYacfmQtYadrOZzNcHhq4SoroUPpbtjC4p5DiClBqh6FsH/wlXCyMJRb6GP+3gtz
BflDvsjz8L0gf3+Qvd8tUmcHSQ8xFVwRK/I4+AE8NfYhDbPUTV2lUJe8x85NNiIJ
APnjuY5XL37lA2BVextFGGgFkE/VLT4Gs71cN9XPhSqCWJnnWUCbLA17ynBpAqs2
i7r8CKWHNTlL3LHq2goXo2DFJbJ8TDi4wQS3whHZ4Xn2fDmLfE3ceBYapw85TrDf
gIFc3hIFZSFPFHnhWBs7NCcbWVaQBoHfhbAyt9H3if3mHjroxepmoFWoUfKb6oGq
r/tJCOMiGL2kjZLWaNzLrGuAA4Umn62xyWqHogOO1di14yVbX1fQEXRS8FkVZ/sR
6nyGKMlxzdIuiYwYlx3DuPpmv/4XZ2aoY5BkghD4xRmR60KtxOyCr/5wWvDNseKa
LDCVximMfrRUrJOjaP6z8AenLB9Y5roULBGw8zyoCj30EAdHqOeHN4ZqFONapKY0
p8/Juz7MjdRm0ogsSoFbTpVgILiVBVp8ZDimelGsvuDO8txeQY29H0Otiz+cDCbc
FyHUOSVo0KXXP3pHuEj5J91LO76sO+cv/VkGOEjJM61WEme1l/8c5mlhAVEk4Uxs
TUtYufBe2focxFnNXxlPQ5JOqeo/2LYxDTNeL7o+Yj3r2Pv6XRMkOddpud6QkMK5
YoKshKYG2lAHoj16CnOsnSpfvudbMWVzA4JoIR/CbTtkxPqqskTNScWPiPZ/q6XH
cjXWELOwEuPBHmSbDdAvUilKJkTa1ZyjAPcxoHZN1h1+4o9UyFX79S1dLx1eRdll
rqGtP1IlouySLEIm3l+kjm6S/mm53rYjY5n+28uE0bJvoDxonxrYIH0MvCwDGrZ7
lNlt0k+iTU/TDl5CrIyGTsKVr8tim5UPsWzmw5oSzhFzbhaSxIpbDdrUmGmcxjgO
Ox99/nO8pXGwVc6zWL+4Fjoeh5Agm7BVxzDBJIiXWhwYKoigcUpA5PkA/Obw3JA2
9KoXzisKhxZSlNbq7yPKK9dCZmx3K8wR0ejZVk7R7B5gcGy3MQjxtiioTjWWHFHL
Qr/+g0bcTK+HsNqa5Cr9ti4LR7E5mYbP7Ae+JEpwUVSh5BX5ai+imCCCVZHDCBT4
sWDNJlTy5fgJfXHuCMEGh6bmsqWudXB+EWQZ26/Fuby1w3jQ3I9ctsdJ7j3pX2M0
RMXqJZFtBgbpunsRHpeI0Lk9K5/78l6nKgrdd5lUuzXndcYe4IM4aRNS/RPA3UVX
Z8Ei415pPIZOLsOE8YrXI1tXQradLDacER0F6EBGBC7+a7mYcXo3vBdWlI8MhGBH
QStlbc5cptbxdMlXkfFb6L3rnGpxq0Nx1B7n8SuERDQMbhI/w0imW9ovMXL3eJS8
zcZGcuIdA1qTg+2sgVAnPHZVNDf/ORguuYpxCg2SPdulF4bL9F5O5B3iCsLcSurn
d8MUif/5Qkf4u+V30FOrhUneLEQot//pNEUhH/CLxRJdQx6afUsQozEhKsvuiP80
8SHM60KoFf9H/ECemOE3eanuLrJbsQXtAcPH0dc7ByrY7LgwWdVvAB0XN75d6xZ6
hfwPm/4UQGn1XHgdCCeE1DRNltGZ+uCyEEIYO9QtmofN/mqAI7VHBuJPyc0xMY4h
kOTZvv80j/lVQKpZkSvknN3HaqluOpLfm/11siWAUzYJEGEjVAnqi+YHtq9zXjsN
KPtjF+F1PWLTBvgUMkEgyCxqg7ypCxRmTKMTZChTyer/T71S5tOy/yrM84bbRNSt
pPZOKDIIr033uI+ZxgyN1sqCk9JH35WdkExnDUs3IKj8vNDu5V9eNpY8sYBsf2bp
P/dHQh5MjB5uMJzLs661fBfAo+CI3AG7S2GGEeUfllUIudukHUiAKZ9JAVOw7hmF
paL/tybJwFgsyE13aP/4rfPzS4fpnB+Q30SOFSzK/4MbRgidzsjbeetatwgYBecs
aFTwTYNS4ZUUeDWUTsX9BBaLweuDTUDGgjonk14Hu1YACGi9fiQhNUDtgXV5AxBJ
8z6y9VZ+KmI9hOPStuG1p4JQswej6jQPc7+nzVf44Bqbm8jfsYz6jvYhBtE+SH4W
SbOXhJw8oAcZ5U4YFYbavCjQ8aWBNplNzfLyLkvcqVymF3/Hh5t+IeIbrw3x9PV+
su6P8UxHDrfU6y7sJEFfZeqdbnXDCLovBGWqWsj2a2x6Zk0Dcxg6DGWKkXwplpcD
8ff1RhK398m74edquI2VBteFo+bOQVsjsqpoCOxZKvfTtmxAWoyCjzbmCUC0WqQ1
H0LrhpQyklFw/p/gIvHS05anAthO3ZHUku6kyF+aQoLi3VbWPc/wSZ4SE06g4ius
I3EnuYnIjlCIkineNwFi2as5hfWUlJnS5j+dMwNUih/OSkpH62TpVimFDatERbwa
IOm2elsHFhq0qhsxnEJ4O2EpyOUWNreakF4S0m200CYl/NJ5miiJ+L9miWK21MKE
H3izqbzh4aLTWY8Md3Yn3iPEDDD0Rh9JjsCKcZy4pTd7ollLleBVqL2WTOh+PuEo
bvc5XdYdl5gnZQ6PWsDbwZdT8QwGnUoDt7HyFfKMXrFMKkf0CPoIboSaOdwfNVok
eXhrw+quGnYNrtpaN/GNckeIZ2SjCcIr7EJ5VY/3uWr3ipm6wJKsX/4Fjoxd+GDU
OchE+t3M6I4dn5Tvjd2cZtF5FqzA4PBCXq9NY75XGGpXYBn9Fbywx7N3EYNywa+P
r6cFzsSE6inoy6zEn9SdbKE9Dfy9ALvvgTj6CRbxo8KDMBhTNmBVIJvEmyIT2dp+
MgyLeWEkdPgfuo5+6HoxXkH/EaHN09puwpQMVMPrw1R7traE0191WkHfl11aTTsG
K5b6SKlJzcTMO8LSJTMH1mUR0X9EDqNR9vmuIW7otf6tThwAFg0l/rI1brLzw598
vRIOgevfgXjmiJD3FLlyBKTaG4iQHPS2pZcuMgx/0iqc4KnZY9+forPuAIEaUXwV
fJjHB7AbQ9ToomKON3/DByI1lNAImGYB809jiQaJFx23Z3mt/QNTTdjjaenMIdf5
hVKOVCG5mIVamXNq8nXGejWPuG83LKqsp+XaMZg7G4FB9SZdlH9Y4eqS+Wy7ld15
pP3/Yx8btqGpwzkL3WmWewy8o81YUoyp657aVR6JxyPJkSlvjtry8BEIIv7pUrBt
j4OvjWREnRy5FOmkwJ6e131nP4P55GVbkR6qO3TfpNfAXe3AsU6fIdPHQPqdahC7
qlMQg8D3JCijPm31aaFTk8RrEHTkRIg21sDY/TIpCS18qkWzQzOtd/cdP2MzaT2A
hByodeRwR0NA5Ne6kI3nBzLlL5OCLO/G5l/SusCgPoSWcu1HFHRYp7b5FSnNYvKE
AYYuMS+9r2C9+I00L2vhokSMXd2lJvdM0u7MJs2+uYQolh6mh21XUccL2aYIUs4b
JYFGCju8wem2qkfEs8Osl8eInPXc0CzAJz4gAHN0YJFxx43fIPpFYOTDq/JEvcfd
Q64MW5Oi7+oVcYnS4wkHdH2aM7LrXvQ/n0PHcloVGbIOl4nPK/zXNi3PsPqXNjpr
ZhSQpZC6gdRaiNph8A+Yjouqte8/w/W1yhEJ1p4r+QgyvoU7G2/4Xbh0dE9Z+WNx
Q8SewPyIN8BxylXGZ7nYz11q8LVkgt1EqGaGzTHYackMII4MKVmmknelAr1R59fo
fmfSe+hQtisZXhXgeEVhD9CSpqlcDV2SOcCoVWYm8RhBrzHkupELNOrtFJLiCbCK
mdR/F+5bhidSukTBGM/qC4V6275GERSd/VSD1FTh2x7Myr1R694AmfCuaplZeWAk
Ymn94pm9Y147wiKXOBX9d+elp/jcOnfzoEQ2wGZLHKDfbCH9BN4RNWCOmQTBbfUd
RXN4q5gfCVG3+e5YHJAtnd/80//RDJA8JIcALlpR5i7zhOD2iQ9rsRyHwbeJPkzC
cbROAVvdWwNHX6KW0UB9KKrcsz8MpRDbbetBSfHceHpx2Q0SPu7vV3N2Gtt04bBX
pXrA3BJbNJhfVnTEX3aSS7NdyQ2yGyEsEDwyEXKj8NSBUdzdCEKjllT3iwC0NmRy
uZJtk/SiUMz68SOq77Y0wdImf9btef1ZCz6lNJEeACwuO5ELc4LfjS7ElC32eLlf
t4U5kW2qdE8ziaXuWcj1WihgyvgIRcMaqI771elVn1dwj6HHnuRW/Ahn1s0jyVEb
O+hNG7Tgnwz+bxxT72oXnF2QHDGTGy71sya63OxJhLJNH/gPFL5rBJdtK/eWbiH+
Wdf2y1NMZ3CqKhsFTXG58dMtVXpwsq3Lg/58YTARxfELu7og859mfFbWxw4uYRV1
sqOJmABJFF1R8nxGn3eUTfxqBsqgMBMrE3fLJr8REXbaXSyNE+s3yPwh1487otzQ
n0Q5JU4Np4fSu+0+i2MtmXCgxYTr0jfprAjl6ey1dKXNzO3ODQhl8WtfaMq6rm/m
HeCmI47pRUmn/879/HqGWATCHtwRWpplzUE9XvXP9klzR2F1sbHcRhSSS/3Gl+Xz
+llPHY0mDpPn9bfzz3tcXtYzZBIEvo3tnbXEqnYyTGXl1olrpaoeZN4JN4zv1UrA
jEESipYRiAxMYilWEhpURKRf1GSS4PCvNfBkIA3JR68J1oh1/27AafVvlCJz8hmz
1ksaXJsy7O7Ufb5afzpNLCbO+ihT8BAlE27HHw0QUXg5xmuHpGf+soh6XmPqLmIW
yFv8MBJVjhqiggPKXrV3W7PE+TtQHITUhVm6KQVorNlulDD07fXVAeJrbuMm/OVa
ERYkx7WYbZ+eQNjO4fRdlF6MQcELjqNP/gJjSOOqfoVZAgco1c7jxjnudKj8AICs
mXMTInKd6SYV96zgVOkcgBa8ThdYxytA3PSyEPn49g0XKD7UDyq7/uZdL8PGAviR
CR0UTdV7zMkME9JiYoCF+waPh+CDUkOyL5rVvSyz9f21ts0uzEdQ6xLL+b+ewG74
LFu7nbxgo+kpLZkfNOnvUDnPlLAyuFOM/INgf5NmRK9xz7Hd0mn2MvsIDoO+ySe9
8E93ZfZ4m/nEiwVdPJd+dpNd3Gr0CtM5FYUyXQcUBVVJ6BPP//mWg6yyxXZzsIuC
XhX0zh/1tPenBu+vbcaxNufSo6iY4QR5fm0H4/t8THsYDzktZH41UCHgT7FQNIJN
OelNfZ+/wpNBGXWiWR8/3u03hHtqCYfkerzwO/vC/0X8XMxHBI1Iuvd8mSylMP71
lHlEWRyfp1oweyzZwtYbw/v52ecToebeKZtwLcgDTBIMGfZPXTpnNAzqiwJ+6tsy
xXs5jk5sNj2wQJJ4dS3VOj4kdbWyLFdfjrxXDQlGrdPT1dVZPPn+TxeuScjPbGN1
MMWBIc/TYvgZ9Nab4W/B/efcECX4SQCHiJBpqYxV5D9XggUOkashMKsf+DToO+v9
wB3wJ3flVVFD0mHW6sVVgLDM36ewHIZnWOd0bOV/cgIm6w8EaYizhePyoAvBNUyu
QOWgZMIZoz31UC06H4FMyOG/GeUop008op4hi8821sZdGfsy61DSKMaBXoNPY7yq
PN0LhA+I8D++jMU9CRBOMu1f4aOXgRRs/eDpfxgiV2C24fmigPbPLDy7IQNhHvn0
JNkCq47tVmBX6fmV3utrs+CAo2M4n8PxdaKTg6JAkrpPwzb2s9JC38izMTWPOxV7
F0CVZFwBQbFGSLG47m8iPfkE5VX2ODVdwPPOLxi6dyltx3OwVEYDOsds3KC6E6Oq
XamuZeMgmVmQ4WBc/tsDtwC+95NaWStGdSAZJBCmYb3G+K8+Wb80yeRlY7eruYHI
SSu9uGKjeXxhU7zzCljRNYRKajsf7tOW+ZrMKdW8N3ye8cas9PZYBCHzvCJQ9GhR
5QoWl0fxgcm5Qf7SqYbf0EtOprnZ+Mf0HpIgIY2Fhk40yzPV75KEYN3Vvq6OVlKb
hlCPXtkq1ePzlnNkUddYllyKOKqLLrxAj57RbsQ61Na7j4pz0BNuhUHn9fH4niSJ
E/d7/F/whyDnV8yBBkDGMuh7rWMS+P4THt/qHro3YlPslG7/45IKjigFtxMFpfjG
hC3i3GhhmjYnyhEYVxNBlo9HkAcTYSuba409EQgsFu17Izo5M4ykQRL83NK1cvsp
5Dop6yyrP9GVtR94rGkaTffon4yJfSsD+4S3cgvODfzK/Yo8HEjqnGQ9HndYRvC0
ZCQ0Mop/44MRhXBcaaeFlwnjEOdg37e1LdskkZhBLJGOJb123e9r3FbSqSP3jUr/
T/h2AzR0w/q4/4uSQxUHHakB7BrmJ+P+Pfo0cA+TfVS+IMERGvPrWUZSlJpsnxQz
2ioszyt9ueLiZP/XZnM8TMbtSed8z9JNYyiC5FHN66/mNhiydZ3w9KkadexX/xrb
H2Fq0K+O4YM+HAerwRlDPQvd88firwtKTfLNUWjcYA9ciEp0VT64DcFHI/gNZg2F
O/XZOIHAY1db+51tJIefa8kCQAlWphAByCHXcXPyFnkFPeFBVIRNBRTWkCUOr5To
8JrP+9aAn2P1XMSwMYaSBGXoQrk7kgQB1PbrmSIVQvv3CE9wbEtwJUBiFjevCcn6
yZkqhxvK3aJnd4n6VnUOfswkARDM6TMAucQ02XEA4siPAekLavCybq1vnxeUGl/w
uxY8nU0s6Gn665WS/sa1utqxK8FNaO0QwIF2TaUBJpXwO1HuL7ZXF0Y5HSI2x+f9
ymVl79iXeyfzh3UjPxasX7ciovxJb0Fgf+B7Ht1jLTXYyyBU5U5+KzAz8vOMIpW+
tE9+W/bQSOc4ZK09cvOSXSkUwqBczwERprSKLt2quIvd9DNAQll89lSxecWksyQW
Mynh4czYDk8ZDeAQNX/s5v77gYLkWeFVD+eN0K+LKKxZHBN5CpbDiWAkwziRMe2/
/roYCsz67TZPs79/rDWp7Ub5p3OM4J0LFh4N9mY13HMDEou4VHIka/sCy49M13oI
r8t2c31g4YZ8AtM6/f60AL0ZmcZo9ZCyWdtGd5z/RMc8mzr1IAjfEV/ORmct3+G7
EQyV6gqOmTmMS/RTotoC22Lq3b8lget49kSVujXPg6D/HFukuN/E2pI5tbGedVYg
gK/bs96m8vpttPWL+WO/PAxydRrSROv+DBjB3YtiKEphq/BVCje8xlquDwXZYvhK
nLLaYyhnUlboJ8ZyvwENut/Q0tVQKavmNh6pwF8k+WnknBbhIGklGwZN5gg9YnyQ
th+chHAEuCdJzSiZWtaUbcaYBcwiwIcK7NELD49COKHkNCmV5Aq8axjQRqxIGSy8
SIfh0TV/Maks8/zQSkF7GxdYrXN7N7z8B0RBOtgkvet64yjR77c8P4XJ14PBqaoI
4h7lG/RE+nVmXRtAqJlotpiGVEt1SyMIesavcWM+rPJVpY93MLdBhSZvaDL7WWbw
Eyvow42cO2y5ZzAEagQslLjTIy5nkXUoUUVKNjx3TgIZvBLE9phkju0iLacKOVsJ
LWYvsMB0KflY5AfJJWzgTPZ1s6R42xoV0MAU4CMJJ1cW8bfhL0SNR/lz5Ruzi7C/
HhL1ZyDDQKtDKPcgxixcdItzeC8mAub1my7s3FANVdnD7qHvjEZnHAfWSvknp4xW
xBCSM1ReZ9CNYqqbg8mdO3ZuP2ypXBv0gFKQsdtIP1URvpQfOmRiqqCCueGgS3wm
RxvIvsKU97bOc3PIWY1IdOHu1lUKMUD0ZcMUfmBg87lzh5eIeZyXIBg6h+70efMc
B+qgnX5hkixJGFNRE7IUxrjbbU7KEEVA78xkBXv1WKAxCjGC7LBO6qP8p3ioOuAr
VSz2TsgKDRkt/USmmzwb2d4EGOiT9PynFrDctDbyBDekaBDZZb0dxGByMuZBXNiB
VmDAKD1Bh0XtCfAH5Y2gXqSO+5vy3btN6oDaAwM0YTpjjgQOvArhlKDc7O4s7jmF
DT+4BoFR90jFIiidq7LKZb+yr6l7IogFmKrwt5fQMVZjKQeYjp7Qd16jRLdZCSr9
+7i+VAt6wfB/TurvtN+f7OYsl7Ezf4weJKPesxIsl7oaQPQNfVx+TIC4l0qmEX7h
lnSUFxYUS8ZovoNuTeQ932QdKPoHaUFORK1rwa6nhX9CEq0y/hVeG8HNwjTmjK57
6ihCDEFaUM6j2VBNiIB6kFH58D1EU7jiwZoPngglI8gcTopd09uzERfpZIV9whfq
b8054rrkKY9loy+X1xanpm1tMqzi6PH//8OKwrxiIeR7zY0t1mUfF3yUd5NvYC5A
j8AcHEVq3/8CWIIot7xyIFzOzeTUhTuqPMXHF5bKZYvsCGB7uqhmKYnzYT5zhH/j
G2pP6s40vhhYT9qkf/PkMtwL6Ro5E/lpSpKwogvCn4cYmQ27Nu+OzZ52bpB7Cc9K
qNMfMk5zjDboOHB4VsMsIkHCyP8rs3RpUS62bqpo4D6NY2d2cne35StWQVX3Y8ay
fu4hJ6JbjxtMLyE6ls423VFHenNqv9y91aVy1xYJnq5GVAtu/5ia3/nqmHWddLgj
2OMKsamwdgiSaUL+HGHp6yWOzJqPCUSq89dl+RgppeP4rZnMdQ3PkFx7DiRgtr25
cXxE0vfREXrHdk/1piZk6ixJTobjntG8Hai7XxJtJ4qToGgInTR1hcWNGghfduMp
WUHK0ri+TkLqgWeziizHXpwForTOfHD06jjvgoWdPhgPa/tc4GL+Osk29h7kIu1t
BnrwiMxAHh26jp4eTyFOJpXBl2r7TTj+em/ZomsvusLjSM/hHOzGHp1tid0l0gYJ
i/pZuXLhoiornv6fCgdgcuoJ+4ERbZ2ck8BH1rS6SUUSBc3N6KnnqMP8wLiklptX
8KQNHDYm351H3tu0E5fTWn4oUUl/PrO3hQ3ya0s4iEApJvH3SUgNcch1GBtut31j
DokzSZbfCrSS49SPt84IWU0pnbKR6IawxuRjVm2vkn/b8z9bC3y1lCFftrNB4mA+
g1qBI4pqE79fJzavqjoBpO2FhGzhgdzX020cwmcPtbsbIIZAAktOzHXBnDjcq6VE
BJx2U8Ran1dse/V3Vc07rgVx4zViqBB4vxS5HOjxi0p9b0t/aZ3a0/l7sP5jM6AY
XL6YALc2J0JbwswOqdfI7Ie2OrwEbUiBFpCm0JvP8Mpp+Nz8Bm9wu9kvDZBTgsWK
P//lDWhx0F6RG9+rTIvUJXnuguvOwY3hiHugetHGClIp9LzuWRza7d4erzDf8/Op
Oiv5ulV/rDLYlgfyt6L32ujz3mSUPEfLVN5SLUtAufsFjxNKTV1KZd2KfM003y41
41MxQh7Tzctgf7dbEYYIhY2FfmRSjJ2UHKk0Iuj1yBwJBiW8BweUR6YYtOePjjZ1
701KhSIsiwjHC8z+xcaV35/53kSUFL24kortJ8N4k6N8j1ulQdYWuLyYEKczPM4z
X9f5WaXaXPC9bKJ0rn5BRbu7LwFS/oAhg/vRJ/m9o0icy02cIGzQzmXgFmSUzFVW
hzOjsNTi9f4Ftsdiscehd8IaUVavRXL0WS/eiwGqvmc/yAdWYSiR87MU74l2NmxV
aZVLZ9gIzX9JvMg5QKJfLa1DSbdvz2X+BHffQKV7P3VpQSykZx3ECSJW7Ch8/eBY
z4NW13iCUEbML3QJ/4DzJh77PE9mLxX3vTSeqfO/I93of2YFdz4bwATl3P4do7Bg
jx2tRFlNOiXrt7ATf0DC1Hr4FV58zezlh3W6B7bYHx5rLz80cPqiqURi9Zmqo8yu
UPna3SQd9ThepVuErJwRu7748WjHfmGnhFoajMupvtuCns1twftHBjUhZj2gCCv5
IRsCB+NkYtlLKXWWpC6egJdxoxQqEVs0bdacRMZFQy9+E6DYgdagHju9enKRqnyZ
0rlaTLZMe6sxR+csLjIUcdMHs3neFT1EmWHm4t2fPT/AEtTxE+bkTxu/USmIAv+1
5wfN4B8bRmLekyd4PkdrxU1msTcu1Rfz1hw0UKPMbSF/pNcpu8BOr0nR5qRGh54H
LPj8Uq3rKkNLKrb3sCmdzHY3IfcLS53KcJvxDmwajkJ/Or9z8n4Brd7w+v5YgL2x
ezx58nZdvaavk783G4HIRuc5pKohb6/vCL4Eg2uimvlJMWrGClU9UzG0Ie9HKGaW
LklvNspxTlN08jBnIJTUDMu+20uruCnpIWl/d5wkZZcc+/jUasMo+/iJfk/cq8Fd
2n8hILAwQo6FZRV8uDMuVv/zqA+eJ2Lc9J1zTzoA3V97UnSmBsK1ivd37tuzUGEs
s1QQ3T/GpvHqX07r8yQ6gjo+j3vClGyJ9bJ93cn5IZ7alRcc6NOQP8R7bcOaiE1Z
tY0Qx13k7MRPEY1pUaeO1n8yjrTaOgIOKsknasBdstu50x25dfTa0dJoXLm17qR/
3HkM3Gn5MdJVsRl3s71Iyu+c0RfYJKVF90uMfPHyuIaXDok16PpmSoUohThClfT8
HvZB1kkvk52n5b+mMkjF20at/vTuYPBTpR4t4+NRsdu5v+h8IfNpMb61BmS3r1EC
+VkZO76k1yoYBC/W7rXVNVj2vxNGw5ITGCre5ROK0PTIhXGomo4aOH2kziC7Oico
m0QZvlExFIcsne4xUnyCLdqy5ijjA9CH91Wj9jmpYe9g9Q1Ie7jigFlnex3WAglF
mOuYd0akGB7WpTe8iGR75itXYqeCiqYOf43OSVeOKHjTmS2eF4DUidcPAKlBfZKp
YvhDea2XQZyyCOS055hNBbQDMrDcDu1PMktxnmKEBPVJ+HNlApM93QE0MDJWnCzJ
PCO5rV2q6CB+wg7np8g5UX4OV8b5oeLdmKsvPH2UIEx6RE+zHjLDLUC6aLj5pXw+
m0+8NOOWBzEO+1H0SU2PriAQqb3VVYvi6EB5ZK4GV156ZrayVFRgaulkCuRVKYQq
1xT98ktduD/vHAPenwnHob8Re1eSxuNCbolRWORwwmF6U6k74/S+kNTf+tnarb9Y
mtaFJCbOez737va9VVViDjk+d3U8028kCgoTx6iLd59/LEdXPQTHy4PDWWKkIpCV
sPt4V+svBuGZnai/lxjk2F15RNnUF5D7APCyNP/OzuStnBwYgf37YV0wKy2G1IIA
zspUKggCSG4qjntZV4YmbvFa+KeNH5jHYi30FLZ5RSiKpJCPKqSBdRRHJmSaMH59
onUvOi8ixSc7x8P2Cdp2CNWLLE2KC/XknrYRGTDUkKcBBijljF6IKVNwLkPmpeLu
tg9GScOAvQuyjlbhXuRXJFP6ZKkDAbfU87ELqbNYhBLRCACjrtSx4ta9gmFyFE9L
nCvKItwgXqS5Nf1sghGflyHm351UoP6Sl6Q6XNlow/1MFuLm0Zmy4eSrZB/tDKW3
kF7E6if7TZhmNqkBRjZ9qaPNP1y+Rwg9qXkge3B179o8sERyLrItuWSW558h0rkP
XVDVd4ucK3jxeVBV87dqkcnf8DeSlOvurFgZSVSzRngNXfMCLO+gM4MQ+w6mxu8K
VHXvsP5LhfbFMPXfw30rdUqNAKY0wTAJP/cVAuyDD6fiOKl9uB5s7634+NGSfVO5
ItisZMGdxTFatyKT2CjjCk8yu1v38Kl3wgTOfTpecCBZ3ymhvGSeKwklZvkrkxsd
c4+8lrtzpvjs3yIWFFno21bNSm+DGQv/f7rT7CcAmJrKQw20132KUqkJwiE6yKpR
L9/BtnTLA7KeiIo4OL3acZwtSzSQMEq5zvPte9/NfUFLRD4viLi2ibhzajrnPkhD
eQde0g1vKof2wun2ZtJPKCCMvbWOn7dCTTFvsz4iPNrv93h7DhHQWIF1UqwnV1KE
6o5yYVNguR2L4DmbfN/yn3eNjQLlTt7YqLXuwkKxMlBYul/8Q/p8HfJMvJYjNWZ8
STASqAh7pYu7+GLUZxJthLtbSaKtLMQJYAInfPcastI=
`protect END_PROTECTED
