`timescale 1ns / 1ns
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company:			
//				
// Engineer:		
//
// Create Date:		
// Design Name:		
// Module Name:		
// Project Name:	
// Target Devices:  
// Tool versions:
// Description:		
//
// Dependencies:
//	 
// 	 
//
// Revision:
//
//
//
//
// Additional Comments:   
//                         
//                         
//                         
//                         
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
module cnn_layer_accel_weight_seq_data_table2 (
    clk         ,
    rst         ,
    rdAddr      ,
    rden        ,
    seq_dout0   ,
    seq_dout1   
);

	//-----------------------------------------------------------------------------------------------------------------------------------------------
	//  Includes
	//-----------------------------------------------------------------------------------------------------------------------------------------------
	`include "math.vh"
    `include "cnn_layer_accel_defs.vh"
 

	//-----------------------------------------------------------------------------------------------------------------------------------------------
	//  Local Parameters
	//-----------------------------------------------------------------------------------------------------------------------------------------------
    localparam C_RDADDR_WIDTH = clog2(`NUM_WHT_SEQ_VALUES);
    
    
	//-----------------------------------------------------------------------------------------------------------------------------------------------
	//  Inputs / Output Ports
	//-----------------------------------------------------------------------------------------------------------------------------------------------    
    input                               clk         ;
    input                               rst         ;
    input       [C_RDADDR_WIDTH - 1:0]  rdAddr      ;
    input                               rden        ;
    output reg  [`WHT_SEQ_WIDTH - 1:0]  seq_dout0   ;
    output reg  [`WHT_SEQ_WIDTH - 1:0]  seq_dout1   ;
  

	//-----------------------------------------------------------------------------------------------------------------------------------------------
	//  Local Variables
	//----------------------------------------------------------------------------------------------------------------------------------------------- 
    reg  [`WHT_SEQ_WIDTH - 1:0]     seq_data0[`NUM_WHT_SEQ_VALUES - 1:0]    ;
    reg  [`WHT_SEQ_WIDTH - 1:0]     seq_data1[`NUM_WHT_SEQ_VALUES - 1:0]    ;
    reg  [C_RDADDR_WIDTH - 1:0]     rdAddr_plus_one                         ;
    wire [C_RDADDR_WIDTH - 1:0]     rdAddress                               ;

    
    // BEGIN logic ----------------------------------------------------------------------------------------------------------------------------------        
    assign rdAddress = (rden) ? rdAddr_plus_one : rdAddr;

    always@(posedge clk) begin
        rdAddr_plus_one     <= rdAddr + 1;
        if(rden) begin
            rdAddr_plus_one <= rdAddr_plus_one + 1;
        end
    end
    
    always@(posedge clk) begin
        if(rst) begin
            seq_data0 <= {7, 8, 9, 0, 1};
            seq_data1 <= {4, 5, 6, 2, 3};
        end else begin
            seq_dout0 <= seq_data0[rdAddress];
            seq_dout1 <= seq_data1[rdAddress];
        end    
    end
    // END logic ------------------------------------------------------------------------------------------------------------------------------------

    
endmodule