`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company:
//
// Engineer:
//
// Create Date:
// Design Name:
// Module Name:
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
//
//
// Revision:
//
//
//
//
// Additional Comments:
//
//
//
//
//
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
module vector_multiply 
#(
	parameter C_OP_WIDTH = 16,
	parameter C_NUM_OPERANDS = 1
(
    clk     			        ,
    rst                         ,
    datain	             		,
	datain_ready				,
    datain_valid				,
	dout						,
	dout_ready					,
	dout_valid
);
    //-----------------------------------------------------------------------------------------------------------------------------------------------
    //  Includes
    //-----------------------------------------------------------------------------------------------------------------------------------------------
    `include "math.vh"


    //-----------------------------------------------------------------------------------------------------------------------------------------------
    //  Local Parameters
    //-----------------------------------------------------------------------------------------------------------------------------------------------
	localparam C_VEC_DATA_WIDTH = C_OP_WIDTH * C_NUM_OPERANDS * 2;
	localparam C_OP_WIDTH		= C_OP_WIDTH * C_NUM_OPERANDS;


    //-----------------------------------------------------------------------------------------------------------------------------------------------
    //  Module Ports
    //-----------------------------------------------------------------------------------------------------------------------------------------------
    input 								clk     		;
    input 								rst             ;
    input 	[C_VEC_DATA_WIDTH - 1:0]	datain          ;    
    output								datain_ready	;    
	input 								datain_valid	;
	output	[	   C_OP_WIDTH - 1:0] 	dout			;
	input								dout_ready		;
	output 								dout_valid		;
	integer								i				;


    //-----------------------------------------------------------------------------------------------------------------------------------------------
    //  Local Variables
    //-----------------------------------------------------------------------------------------------------------------------------------------------
	logic [C_OP_WIDTH - 1:0] operand0;
	logic [C_OP_WIDTH - 1:0] operand1;
	
	
	// BEGIN logic ----------------------------------------------------------------------------------------------------------------------------------
	assign operand0 = datain[C_OP_WIDTH - 1:0];
	assign operand1 = datain[((C_OP_WIDTH * 2) - 1):C_OP_WIDTH];
	
	always@(posedge clk) begin
		dout_valid <= 0;
		if(op0_datain_valid && op1_dout_valid) begin
			for(i = 0; i < C_NUM_OPERANDS; i = i + 1) begin
				dout[i] 	<= operand0[i] * operand1[i];
				dout_valid 	<= 1;
			end
		end
	end
    // END logic ------------------------------------------------------------------------------------------------------------------------------------


    // DEBUG ----------------------------------------------------------------------------------------------------------------------------------------
    // DEBUG ----------------------------------------------------------------------------------------------------------------------------------------
endmodule
