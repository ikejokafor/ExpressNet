`ifndef __CNN_LAYER_ACCEL_VERIF_DEFS__
`define __CNN_LAYER_ACCEL_VERIF_DEFS__





`endif