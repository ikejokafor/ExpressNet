`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
62hNKvSJThPlnuSUKh8ydmsP+mn63NQM53CptZjvRUq7Mx++LqN2HAQJVG04Tmvp
uUXRotGedrpKFqbltuFip4Pp/02TD9KtwnOsaQf+/hoKnvsVPPIsBZq4as0znaHF
XntuyeXwswXqCGeg7wEpgjBM+QRf/LUyG1PCLqNx7zd1fovKtgC7UBzLHd/OXgkS
IrvAaqewMqBQNUdh+pFKweifDQ8Owt5NtwdwoZHMS0ACc0sPAWyG/qxFoR/RUu6a
18uKpLE/64LN/BYrqKCQDmJxV0ageDxDuQwbZm3GIvJsV+B1wdAxmvRS08K50LrS
MRxYgX941b4G2EexRE5ND5NO39W9NOgpFczi46lKYveFXKY3W47I+jxL1IKcotnG
dtQyYF/o5NgXyUv3hZeqTbqaX/FUhzrSxN3O+HqarIfbvqR2CPJh28X8nCdVa2zM
MRO31XPDKNDXUu2IHlzgxMRh3zdF6cXhB1i/M5pC11QaQjZjNvC2PQZAso4VAUw8
iHyG+A3mqWZZnr1Qz7mGQD9nxDUGMj51XTn0D7lUAian/+9YkvpxZN4Hziqih2gz
diwCS5OAQbKddG3OkIkIiRTewDPI+ybZf79ICXNj8PpZPKP0vOFhAuTzWhu+HhGA
eQ6Z9s98Ru5lsLnf1sHSVP8WNXkh4WR9E3TGrFt0rEI/XPRjsI/DEi3/Y0UeiHSh
iA9KI0Kwqj/gHY6LmKMRpi15uRLhTte3q4eCER2oIQad38fkHuN8EuP+2gfk1DfT
GrJZ/VZ7sYx/ElPG4OW3PUiwM+e32mb81XTsausN2BUC0gcXLH8Xjsw7YJA0dbz9
rGwNNDAroKGjS/vakDhl/QB0OC0//VJQqg6nBg0FqblI9LZlmd0qHqMjM5ikfc+W
BSHxxkioFixLkapwMe+syoEW0fKcrit49zfD+loUcEoAMeWvuoqMeqsyu2v5x2AI
F3IHR4fEeDhwmiotm4IsXv7tB33U7YE39zWMBi9SZK6po9+LvfofAocMEyVKPlBf
GdVNjIopEPAl8LwNZr7byRJChutroO2VCm/BJJGFMY/PYCxpZGsQzhbWhm5LkGwr
whNngKI8AHACRbXFnXvqbQEK58wBlzFa/j1mEAVaF714lM/E9I+dMh8LFhnCZuuw
jRu9d1eWVdDnkhq6RzJrLtOHPfTQM1PkUrG+UgGrF2FVDEoa55Hh6VZA2OuUhbds
Lu9VaS0jpHHm8gegQ172MkdeJGVrvcmNjmtwSac1+9Ex3AX+ub3H/+yiLv9TBXNt
E6XRlUQju9MdbCmSF0hI3n4vDc0aq2dkUXxZGV/KAIt8O5ZNrNsfv3B1uF2fpuJc
DE+l7iF77wiiLvZ02dNEbA0SJhGrTImvi1qPgzbIg52EhQJCneKOU8UXEljsiHME
GzA6PzGwUKcfUsnmzKLQfD0ahgPWeLdn84FyDYmF/2WXE6LGpUpLA8NRFgfHj+Gd
jSqkg97CjaEjlxX46EHB3ZK5d7SBqWBoMu0JE2aE/NOcfgmUUR8e8Q/ycZZ4mhjk
ni3/zXwCSaWpK7d6xlXEFgw+92m2Uf7OoIpM83CeccUEp910kmBcnW5shWQsByPY
dnJZKxZmzAV3knNusKL7rGL7LDkccDkJ18W8vQLITweZ2M5WpKdKzti7KURP6pR4
RkTPF3Gcpyvfd2DQ0DzSWA8lQQF5cqyYSh55/gBRNcXelLK50+4z4s1yR9DMvi0d
73w7DhQC3uMU28BAlBDxelWs5kGJ7AnIR9vDOgrohFe31uAX2zvLiHbBxydfjRNy
rjfsCVS62Th7lWia9FTEm6lfxfCKkBgkF/sr4PeSiHo1NO5WvURuTG0aUtbRUbdN
s0nfh8cXy9BU8VcQz+CACQrk9OH7Vzxwrm70eJHChMamIJAL1ktEn/kf1Y0isMhy
pZN4uDMWdLQ/VbhGgrToMTbZF7go9f4Tz9ERNdRpCJItKiRS59/29wQjgpaIa5Lw
ebIaPdfgUbFnhezrFAZcd/SVexLQr/dZ/M5nrrLiOsZ4aieyoKSzZnFlx+PgLHpk
gXhZbnwOUzfKsuHr4+9M6LTT2QGwzPPxZ+3vo5ll+BAiOwTzQNTNsEOnXERYC3s3
/IUG+0UmuTZXtrWYYYxjqUk9rlr35yjcZg7qax5n8enWzkqgZpxSijXMAlpLod1P
WpK5lweQ1DDPGc8Pw9Q4nxDs7JbTSTxDXePn08iZKtGOJx12oeokEk/Oj73qL/zX
DgLKAqtNXnQgm6nvsCbSp2uN+XpHwpG3iECiuG58sMgnnBUHzQvc7LfcFA0XkqGx
6U1/aYkOZUHwxeBSJlH8++YvuP/brq4hirppmUc3JRH5Qtxdqhv8nsDPRF5stQKl
g2psYdgCWbxmFY9wV5f3dXaYayIFwRMO42b00sjOXM0M8q6DST6V2X6s5xZI/tnq
cC57Q/jyB8s0j3O1rWyEEVWYc+pmFPkIiIumuFZgj99D9Jk+Va2lz4lwTSmc3T1o
TsVx31rA9xGAHmER5HLYFNkxvCcyxLgnz++iWHv0ZvMdhRBYYkNW8qzKNk+wOJ3T
w+4/IQshKU3LJ6vP1Ei+9iDbUraw00mljVGn2VmFN8SEvL2zz4L0jPCg7FljoFAu
cH7Q3f2o0AkKJOrL6XToVxn7e5LVp0v9vxtqNqe7zGpX1sT1qPnD+CObVhAwT1U8
n/grDcyk5PFQcKT9Sz2UITW/TLXg3wP4P/Mss6Cl5ZiNSskFqCWJxNuIySNt5waM
VVKTB1jPOEq01SFmC5z9OrrpeNAM6eppjWhhz+Beb+F8660UVBKOYgoh8a5lTCN3
R4IIRbEm2W4fB8qHFn8kvmWGpRuZeFMiYiwtT464fduQffSYENVnY7ODmBF1JmPh
fqOksNlw9AUDKRIddX3916BHiN+s/u4sWpv+nMzQLmO2GmFbdo+ZTT4898/nTYQF
3lo08PLU34QeKi/GsgsNgRM+/qb7yUdhrSrWj3Hr1EM+nDfgOiyZ81ZMpo+oJBF/
el1/gYhthfLAdLh7hAnAN/qMxeCrsvYzuYqtNGyt2GgZ0MPWcelgYd4f6L5pzOS8
UiPzZPqN0buTEjbNu0aMHoAyGQAfZGMtfO7DbBfBkGQgEMDOzm/HhdJLZc8Ig0P2
O/cYumcBvjTKC4u6DJiQ3sEnDN2h5LbGke48tMHvvkyVbXzPDq/ikhOHAlbEUHSs
uXmcp0OS9epluakmQQDDJ3Q9S40yXiPB4TfSSyOUA2x6E8ZfRbTnwg1A7xqksbVW
a8KC7WhU/OeKVqJPLPkoP0ldYxOstnja0Ln2U2NzTuPlh0GDOQUUCvAG9NU/xEvI
L1ljhFJCBcAdd/S2yuSgd8RF4D11SU8TcQKmzOOR8ZTBNq3OFE94zQ+/5s3CyOdm
juR0HhBjINWIsd74pGMVN8/au2Oiy/SkTDBImL4pyhAO263I//FYKq/VT+tQmvTa
9sOmSKqGc5dEB4VKpDZI8ujpo52JjRveM++NaqftuSyhOzbiW28nbOWuS2Tpgf+3
lGuuY1KufEfRD8/T7OJGZvxF22/x/paTWiigjTsFZti02bDFh0s4fl67WOsdtp82
79NBqK0yu7raWUpw0Rt6w1p17XbqhiMPayy144I1uL/lAvjdgZXzHVQeLKFi5xtP
FOc72OyftV9xUaKMw1ljV40PU7Ux5z4QneYSigiWSHEmkSqdRegGcIoQPPCw0sPj
QQv8zcR5hlbSxcg8G3tp1kzXvY2huPCTecleCScO2rbRw8iKDRDZnIrsAzd/JUlZ
gdzY/yEERy2guLfBtSm185FhSnPQuGc8hw7I6mHmiseu57LqSB5NpPFq02BvX8zA
5NAKOMCeS7guZhG1MspR9AOnhw7ne9z3DrK0m2+p5P/JFnHutYkI3FmNR6KxzEzI
y53iXJpDmgUZ7IBUWOclBBm49suVwib5xs6xdmjtUHxdqkibEhc5DRtmLLlwjAYk
oH3hjrFNDs/L/nG30upEWZ+1I/qmIGmgxPXFGkYj/EO85CRkOfhVvGsmVTyTAFMJ
824ySiX1c5Vef21XjJMz6BNpG+pKek5y3BZY58DUPGyQ5WjGNNme5p2gA35sgX38
OCRq+7JOrhBxy8ZOb3RxuZiO5pwhCTv0VJXdHEG0oRxCykJp6QX0VzlmKDFBleHS
lKRLX8oP90lYbIMes+SEQ5P0lHaCVESql9ihPIZsdEanQOEvo3E4Tlg34/B9s70m
QLNwj1AuRa6AjYP/2XU+GUmdM6OecII7DOXXO0EH1SKD/rspwW9yd6uqCdCHt80A
mmfXxiD9qGGFzlIlHfNiMhphEKlID5uBRLWen1jYm4uf0nvf8wUs4EAl5c1NXIg/
I1FjFPRkVjeLCGaEI1n6Yp+vaQH0O7PGlyphouL7lkJWgmEwF+kx1+w6o+TeWlQ3
dYwE2fUJKbOgC+/jlr+YnI93pSh1+PwD5rFo6abbBb7uAUkyCPlz5A/ID5zL9HZr
U+za3GyqNpbFm3m0gGxNQaTS+CnqPliJVO5+DBkEGZ/tV5AR0CT9hMnPje/FW2I8
SaMVNnOl1SnDy6n/0rcFcbfFrTJhdEa5rv98vk7urSfrq53Xt4cgVwgaDjPvdkCd
WQKWTZXAqhjLHUL71pdaTAkkJ+VEEs3X8ow3hjpYL32N40NfLe+ubXTCqgoGOlgD
n7XFlJu3DEimnI98yFfSZBKTzSmOn4qwFAuOLqonQiwRLqjsKfB9hdTEO1lgcV5N
0sg43WFkQizOu5jy3nH7865QI3HHJFEvj7Cht+lpnvolotyItX0u47QydBrDZEBm
Zx4cZv5c5cHyUQ/tIBFH3EsWBIyOXVP0hfgSJqNqgqgARPUXqbr6EedVP7w7KUTC
Y8y85YvlSUjAOEMXHe8ZqfF+06pQjSxKMO/6qljdWoKuXP9EklHegOGSWtGw/5t4
kGHgvNDyRYBS0eANF3gwxWI087vEx0eez4MXpnZEu5vFCWZkbZSdQrL08RxgyuZk
F2IDlqEMVrdbeDlewBv9tV15wd2KMRY7UVMgUmohHF0uwcxYZniiG5lNnU3ChQFm
ecXPov5l4yNfmcJ2mnCI8aAgnZ+PPcyVDIOd2hP2DXV+MKUgyxn3XCVi+XBWKFA6
LK1DyaJZBCD8DpOnIcbk8vCtHEIIJ/j7LLpoo+xjEHJ2cOTZJSkTV1p8ZoeKLMYs
mk00SA6W7ebU435tutUEp4Y7KfMh0kffJdngomanXp8Bt2xv6iUCTWz7FlYJxN9p
EM85SpZOf6KXs6TmpbvjjTpopPbEB1bckHPHXBy9hEOjpGWOqSESBpKPzurCva3m
gpkn7eQNJugK+nwcMGYvTUaGJuEt5hlaZEi6M6xKk/hi8cnOC2GyAIuiWK8o2OhT
gJ2rftXDj2zRTrXr79S7vyByZi/UyuMq1V0aLMk/3Q6I6rEwKQjQfBvQ3hRqqZAv
id4ewLJ1qQ8flkbcFDIK701Uf7/wzaQqa33uJDVkTlKK2UojoguWTBkrrdx4S+OP
PWQcgP3qvXlappigAyl5HIeQByzeykU6SjrU9kLejn3lObg7IifLGNvzn7hUx/Fd
rTs1qBM3a+kiJ1SzPHitWKPK54+ctwgsNsOSC6UXaHxp/TzuAXwsv/QGWzvTDHqj
wORYBIzECLcEV2nxlInlh6KeYoK76Q8IQjmmyuePxtLSfeTiTjI/Us0fFdWhmj0h
EEUNW9/uPYHRAqVVwaRO3+FKcDeHiMpNkpd11SXTTT/lsxRFsHLB8/NdZX4YCUf/
iWSlKMQwekJlpojA6UchjEwcU3Ncgv2MN/C3bS3JTPv9XeANmvx9AqIfC9RNgwOb
mQ4rKLybzniG/BN/3i4RBkIrmZ8dV1jRKIwdEPrTco8BdsBhxb9F7YyCmkFPku5+
5uLtqNqCPY4gz2YJvcct/hCJCtGEm/oFqV4zRApE8chHeADWj+yUrNoB0LagX+BX
uKc0iWXyGkwMTHqme1lEwIGGHFm16VVVJ1ZvCPC573rwJTd2CO9um48YsOHsHKGT
iJp5vgMJN1/opjhvudPLe01aDBAQhIzQIE8fjpY2DsZbwHzmBDZKpGz8YrmZODCD
M0HUoEVtzvZQoCGn1O48JvUhDec/ajNIN7OOVEeZMleZ4ccOW6AxQhy2d3aR0jZE
4NpGL0KC8McTvAaaprOAp/rOKn5r+0zg5dn0QoJ1lDvmAkvHm4pc5Cf8Z9Jj1851
D+BjaBpTC6H/hPDnSepdy++8PCRgJegyNq/2sYV1uRHEGGYhHOLRpTqh4GTLQ1KL
jyPfcz3FLGikIV0byoYm4vykc306dJfYI+ne4YqB2555S/WHAk2bMdqLnIsF8w3x
D9cOiPoCEB9IzXb3i//6q1I7wTB0TubSm48ixRx3UlYjci3RsiteMd/jqm4Q1pzS
bCpGqaBvlfyizYQJ3f0amMlJRCLrDAfJyk5QeiNHaNv+P+TmNiL7PZP+XDGOJu+u
3VE2UygKwsd4sksErpqg0E38aOl/TizMM7ufr46xsJ7ZyYetZyoO6o8FZgK0b/9E
xZ/nocqCEGZOXKTDQT1PJ4XffjxIq2BL73QXKezSsmeortOhNM41twNZC5Lr0stv
XnYXDeFNKexYfazncdm6b+uWcpa/wMIvhJMC67YYF4z19j7dwWB3ATQsahaEAwd8
wUo8afsTA78QM08isG/qAyK+YXkFaxyKkoLZqhUyw8o6G337u+BlIwWdcaidymVP
RwLtF71RnT6Mt5Fop5kH9iGUzPM50ldlvdHzIhBl76dMJui3JL1xMzGtMNSrdT99
QiTbz4o+t4QzF9pQfrgs0Cq9quv/ycidSOStYTyiuGDVftFjWj+M17W+P2zsQcfY
b3j9rt+Y+yMzDEdtGjIbalsA9vRRmIffw5528Ir/Q/INflmkh0r38+AhRmwb+fVX
BcrzW87NTf0WheAwh2pQZFFqG6g12VdaU7pozAN8doVE/gsAjBdqMSNp96IkKwBv
19rdcnx/M+md+Sd4eo+82s1w09MJ65zasRBBc382BKYxfMMi8ijByu6ma37DFzkq
v7+nhO0ljUYUGn5kPMfNu/MJ5epe+B0JLqogGdYv0p/1+tGoZp8zEOg9opOmPwIV
5YNppAR0p4IlLKG3oq8r3vdSCElkfrNl1Qi9V7bZe6jCX9O0es3SinmFSKXz9zaO
dpi4qH04hjyaFCcTRvHMSnDyUEPjjnOHvKFc8CLanJm3b2MyKtdfSr8+Jh/5Ye+Q
YbaVrLLjm33lmgzT3AsLYWl+yYR8qq05/yu8iWb3pfHL7IhFcRZ31WfxOhWIzIUv
NdU5OFcI9eD3kY+JI+YO6MJCafY+kwQm9OMdFDH6ZwzHkkaJlLK1fnyuTIZ7VGpz
3ycodgSvi64xIuUdcmMxQGEm7ebEwrlihgRvKxnL8cAkLabW83TTHCz8DxQAWR4U
7W0+oGdgrsxP8Qx2Tet0wxQhVehfKURvGtbdpXGPCPlKqGdy19/uCU4m3TD2ynRN
nXhMZ+vB6Qvro88mXWSkjqDD02RLPGjbq6t98jAMK2UkUZ45FR8XSYJEaIzSGXCC
nw4g4SApzhcMqgA1wntLsKDPoPdLrfjE5OVxlChrPzdyilZNNq65A0fTMDlUiVov
nC3KxdLvjdMJq1EJgZ0CJpIhPwgB0Uv+gLx1slY5kgRmHv96O0/+wL78zKpCUM+s
MbxIK1TcxdTR1qamx7TLcqpiFnZfLX5Kyrz3gXQNxdB4auzzGdb8mHHaf8DN7tVJ
VGZWmZ6EC8X47U5ysrlMFDLY6ppn+vEOJEqdaUx99wzaMuOmwsVaJz47wPUj7XQi
eyyfgoziwqB3z9Hksb8a2quK41x+W+hBaGc1azUuoE8YbtS3aiYAhkegDlPi8A1g
QjJ1KlU6yY7NMtkRRWYCQmUhQmN917a3XZCvEGHB1mrJblGjm1OZQ9iKNFUJiBJu
jQGgtTz2XMEX3QOFuVDsVjICAxqT1XSBPL7RlY9iBxvIG0+7EKrHQ1msmAEdtBCv
loitu/1aRHzt8/PjFz9VlxY9N2Z6NDOhpmalYV7+CUOKMgTuiNG9m0jmmZ8KwSWT
QEAMRkZSV4XIWEGQVcivOL217BirsO0cjV4sd4yX0LaCNGYKaY7DzVJApXTyaChU
QDhLyKrnCpw8IKPLBiMLrsxf0TYCq2oAmdlvabRT+N8yv//JyXEOPWzffZY9MZr9
NI73tuimunmmP9poT/ltX4y56I3eEA71AfvwoeFtcx2OJ9qpjvKSmTrPo6TK5/iC
Md9CF//paKYFq2McRLaOhsZyHVMOSL1WDNEjaoK0Mngd5RBv53u4fi9Ndjd4LW9b
QjC6HNyS64sfzQumDvphTvG1IMF1EOPq8Riyhn7kANJTGieoL6o+Q+Hx+CObuvCi
DJ/XL8VkL+8uDgc+x4k5wA54l2jV57j2B1Y+hbG+wHUH1674LCJY+5CgNyle00Zr
TrRV521Nu5eMkrnNS4ELsOoBHkJ6tPHFFIl5c1plXC79ZViJenWZVVd06Qo9jHIQ
gbrluscjRe9yjET6LBdYvrhfY47IsY77JolMJhY95riIItGNAX+sUhlK3Q4sP/rs
2rHhrGVpL+2OckPB0rWbsPnsC0Esu0Xl+m4qeTDJvh54VhsXiK36KmCkvdsGduLd
il4uoqAwQx0AFkeMGlxd0xdUjnKvX7YXdMCpy3imEUJ7t6I6wEc3+y8nQEbwDd29
2hVLgzyJiYIXzWkZq6NMv3DI1jzLwNjdNybT9rylduUGLUvrnKwKfNfwwyQaY2DJ
m3u+QzNPnQZ2zILkwve0/3svfq2tSF1wtZsS/igj88uAR2ZThxEKJ5BiQDSdJ8sy
bDN+IjNQVhCqSl5SlcTLk34d6s6qLrScah6aZbkdHl9gh39KcX7BnyElYL/LvjXA
gyEBZxGttO/u2JMYHFkMS9EeDFtzXAo2MjFiyE6PgXrhT6VPg8yCOEQRjt7dzNGW
Ceo3vR2i5MrpV28ETuVIpJUZ7UTU5jC+3iTGhiuNZvAZRVgQUtojXMEEHnNhv8IY
yECp2b5xzH3FZ3leTA3sAk+DQ79TqJS+NAMnDN5bjPc3drJo6PbBjFUB7SWkBp7z
5lmrTZnYtG2PeffzrFmLjuI2AiIq+0CrBtZdO4ce0fY8b9Zm+FqFcDgy+IViEi3+
0669BNcktublR8DRuOS/GUhhaI+s1DohrV2pBvG6tBAPqffS//FW2bf6CG+zYiJq
OErPJw5AozNv2Ku9XKzx/cTxzXhCacezw5iHyOXe7cnTqSE1HfGDM5H6mKK6RM3q
vhAh6WpzTOwRgrSmj2n3Z6Kk9NRn82+rf5PhCHJWvH1b8+FZo8omPFhIy8ejfQ1j
Fi/rP8qPQqQQu/lBAsaDz8Wy2HkqdwMh8+tCt5pvEucTiDzcWolyfI7zwcxigW3C
a54D7SmYty0smtkjkv9S4M0DAMPUdvwT7s8s37dJXh03Ur0z3jt27A6UmTStCjjQ
G87vzIjfuuLTME5F280uvUp18EbS2knVgTAy+uGEN+4YXYzZXfJniTCqDNHjI9ie
Zc2UqTR1ZsTZuN6ohQ25Ko2lrYDuU5BFigCG9Fq/L3Gso9ZXv1xPrif4ZFSgepPb
tKfRramIDId3Z1MIAIHNKAvU7z41p9qLqZ+GAFLvJXsUE+8bJDbT2n9EfZ8VzcnN
trXzNvC8KZyOfYeN+IuFrQzmVAIl0ILJUKJTW0qu1yWQbgpCEHeUpCUmTUHlRAnp
9YHDBQMVfN6kPDAS/WyFdmw6Ooqd+rmcijTjkOqP89UabXpNHR3DIUadI37efZuW
jIvkBGP208S2dgHU4vCbHhZ/MK559PwCHbqcymxpycey3L72nmT5jhbtRUOaXqi7
YHtQif/NM+O/QWpspUSMui7VxtsKbziXKvQ5BJvsvsBEs0cpAFRlHDxUPoIkQXcP
aZTmyl99YcZaO8C/5No7n2vmUxjJsMUFkyhuyQ/xm7oFFSic8ph2tMLnkQjAR+l1
QP4uCb2aA1EIx949ALZRoSrUIcfeM5BfI/RxMDKFjL+XFKfRMEHE62VKCkp0cDE+
6TpJ5njXlcWoijhoZgYZ/xmscHbUsy55UEZ/b0RerDxHWt6KBj7RhCWFYZtQhF4E
rqqRwWSPT6PcsvvvtrxOb/dNTswWC1RQ25Mj2eOVulX8PldutLmnXvUqzUXYHrig
WQB6DD1V2Jc+c/+zDDdTuVrBYVAmLD/FPycCJs0IVbM4EanEcjTR+q6SwTjgMve4
c2W72rHVwEEWigq5DOWtsBj7UTTPIHBKMEhdU5rR/r70CifNpJEw8MdtacRzBOLe
uZcOUNDM//925uVjW8Kynu6yTjDTGPWBN7jvNmLPxSEj9Ug6GapGH8mjmB+VueXI
/0FK/hQdZCfKGuP9RV11hhaBtvw/qsHYu/FuY0544ZfFY6REBFgO/NeTNIox3zbo
876dWX74FyCSfZInQMeA7dMPrP1HXEKZq8uWJbREbagDoj9rPtRZDPr5iBl+itbM
i6h34IQMUD9wYncIBLm7iSZjWYicSMnM/4W85f8vhMPIYGBBxwrLgOneKy6cxHZI
YCJlWok7LWrS8xI7lf+4Ce61kZc4WenOSo5ujm5qPnV3CR4BCBge0i7pzIdCR487
1Ds7sx3yCsUxFgse9+h735AZQt2aYIsVehI1Y2znq8p2RAvMRrm4iMLqNV5LIzAW
fSum2F5pHPg9Dw7CY6BuPnoavbV1NYozBCvI27uRwvw7/uQ0oiZdEhL5pSzyobOB
ioSUU6n1Ef4xzW4AaqK3AXk1+xf4wPjc2Ka/AyRr7Xt1PaTn+bHllYIQRPy628Uo
V6H+8tok+k3+4fsIBVNDNLmUmyo3/YXyG8RuUSCD86qvNdpZKBxYy6g1x6qwfVWk
YSXjVf8ABwlUa/KCGlMoLkwL0sHbjJIwFwkydUJCb2L08sl7wIObX3bnbWXF8e7W
8yl5CE9ZXN8+P/pQK3juj1OS+k6BEwFk4CfCcPwxIw8xURBKLBZwk4V+Envb/Bzr
8J+0Uo0KAvzTpGUnPq88wsnJv614bQhFhpbJj0jgnEguYPHqsM2txV2MiVB/9hsQ
pAtFHri83cDF7OfzCuUgUU3vUherMlQA/ELcv4ftgiUTA01JdHAUkaDjzixjzCcw
MHCBD1LXNSXWgkI+FJA6SQ5so7OFA3b3X6ZdKyW9+SlrozDmxd/3+FwSVy8z3sKg
7x7RouacmYy8xqVk12XR1ONvofmWH3aZtV7QGZ908FIf2Oc6bMkvHRHFAoU3tXq/
0Bbc8qHBCq2CsGfYXCagStguIUXJK3DxNMZlZXXkCc3HeGZgFUeuSTzk8PqEvcIw
N0FRpw9+riS4DPGMDNwbsA41JK5ehT+2y3P52rrS1wJAIRycgJ93Psnopw5yNr3n
p1PwgOCV7wEQuW7PE1vlRhR5IR7+1IUC2VvxLRQRf0/0BjQnsISvJVS2fJ26Pinn
gHKYDOeQqikM0w2oe3qEbPfBZJQZE1YbvgKAgPIK8pco7yefQ8+EwFDgn+8oyvy5
jQwqfLvLXdlWfZ+RyAuCH6lkH2fQHeiaIt6yxKoSmx8eAtGBqP9B4zINyfubP+jP
152I+pGQlYTevZvP6+Tti5puH/5D1++qcX09f6aE8lE2IsXVJNJ4FNQBX+w5oOUe
hA/mDpKXnzABogkscdx/qhIh6E6KLD1QvFeX85j6AAoYPbDTHoe42CRuNoa7F/3S
ravQL+19KektTE70AxD18bGZ9NQMIXootcp16j9VfPn9lTeeDqnL0mZATW1wTxE3
yZPmPOyx6BzYL2wAIasw7Z8hbp3WWM7vcs6HbwiFivgMceFhyR4jQVgWmdu35Fmf
Gnt1p493yaZLP+R0YoyEfgl6TXpkanEKc6cUqukGqFo9gcfo+BRLn/udcF9ydaMA
ifEc4oW7k6YykPKfECjKuMI/4U1eU899ygjIeskIpckMIuuq2rb02JqdpvLwW8/o
HzCbP0I51KpDLaZj8J6v3s/h2z+kq8vvo9TQqUAMClNIK4dvMBQatKDt8KNXE3EG
H++4UOW79JWEJQRsT+dWQL8smd7onn4o8/ZwvdUzhV1TIjCfIbHymgnlByizssVw
5TCpKnKCee0sR7LQ1BYxs2Go1+Mh2X3eBGmu+/V/TXCsbLRKijYgbsXlcsbscv8M
zHHGe4fvDTv9XDof0L6N20k1xXN0i0GhxBxmLEUWvZcflk8UdMSSjXPL6fyL7ig+
5EG4Ntcat0M7UkDHhYfve02bgoBqimIpN3gZvykRv9h4O0lGuRstUmQCAIsfBU3Q
2e/B+a92O+vZtkd3uMsMGOmUgez8hlsWYlbHI9Fuuh+5m830LhWRYTZkOIu7MhWb
ECT5Gxr2GCasyLQUrOCmYTrnTFlRU4MSoDkUWPSasT1YgAOfhDniSAuFHMWy6fRG
a/o6B4I6RMffqAr6XUv07kqozu7dfI5XvHt2Ey/cD2ymTMH9pRvlTAI9qjOoR1jf
aWr9NYIUMX8kT8z/nCltTTe1y9URqgeVoKDcx8yfaFxCGRMUsf8kUB6fekUil0SV
Du3MMKf1fcpZhnV3dVAzkhp+G08TZDInq4UItEd/TpfoYHCUabZ1BIzRA96+HW7s
oW0wytvl2Acc2U1x7wl0dJLMqt2lKrkW4l6c9yxMngj5qYy1gZZWq2p/jb5Pv2eb
tUESyqzKkf9iVgqsXUgkcprky/JcuiNKunlOwHGayFpL4IwGOBJO3zhhdA9ki7TK
RwcbAxQmBJP8C7EIeofwsLP0Suikg+tkrAFItj2Q7S32AhOUMxBrkFEXgxSXpAea
ATvm6CX7LT4dPxNB4XwmigM242LjT7XffwNZC//iOKIx0V/1AJqDMNtdNhGsUFCX
CeNeIg/aCZsuGPS/QObXQAJn0L/zHIKInj9yyspj934Y/gjeUjV2Mp6MosGAYhmq
Lq14XM771t3/o8metRafZEH35YbIQHTT83T3zdoaCsmEahup/sEvIc1bDh+zjfLi
ucvSlpMYU87GT99ElWRO845v3MA+LwE7y1ep/+XZW536jA8jPBPoeOo8VV+8SkjO
BPYeqVF/rSLbuzeuvGntEM9P1BSeR/5/qaaqpXzRcm7h1fVYIqP5qgW7HIFQh32/
paJA1XqvnuwLxvk25iXoVL0gUlB1fb/+sDSP7EpymedaLyTQUdtnTrote78PBNn7
AdPaVmWvPWhXl+VRMEbhbmpgx1NyLY3ZP6m6y3nIcPgOLdMazRkiXAHJIvMaeT7T
wfsS7tNr3Q3d+j5saZ6iiFnZP4i9VoWJksJY0CNTZeZmqWWCvxzTAByJ4qlBVFr/
f0nTe5Ot2NBSPtRoqQxSFFLdzY67A8LsYlnpyxpFIkTwMA0jHKW/G2sBSuGRkZg1
YRCsFFsN9Lme0P0Ok+hbS5Ij/YtGr+4r2N+96NqU/ZfgUNS5m1I1LexijwcwNuxf
PmdoO9UT6GVel/NYtSUw7S/pDWCYK89JFEk2hGSm2F3m53oeeC/0FXfHo+RWRmdJ
IiZOmoYrO/UOTEaDX+O/3lfmcFQwpezYDxvXG/gcC5djZb55TvLM9Q3aC+Zb+nW3
PuJtKyMRP+CacQee/L1wuypn7t8CWnuRuTobj0j7sTW9ethh3WrJguOHAkvKJAUi
eTT/54ksYVSOs37EyQ+iRWzxzLF4D+8eG6dKmXt7zi46RtktJSNc8AW9sSzxrjUR
BPotyp1bWbNyZhgDIwx+xV+JEXMp9Oy9s3ERNNCQOClhqL8k1FwdLYevO4xWDixJ
4py26UFxl5gDQUd2vg+TVhu2iZrUlgqizItArNj07ySIbgzr+Riuvqb0UHbttHLI
NOp+kLOQKXJvzKthTOGR3ZOSpsgX3bHWBzGK0HrxtIFiV6+iYV+yEnn0mv0tecN7
OZ6wIfmoXYAfaAh5ebCWhmAJgULAxLozKjEjdDylp/0dKzoPh36RCNz7BBnc0LUw
2f4dKc79popPeEana3BjGoVqgQa3GwneFrxBfHbpdVpFtjFlMo7G255XQYU4FOf6
jpDNh8X70cgQinLeyd6WFVTWBSmhfoYQlzxmFJp0fzTASJI82l0ChLN8mZ6qG9+K
E6OIDDZhRm+KiGSd70zcs51rLIiJ3OBsejCHLKWLEpFbylFCPTqbeAktqE3hzwAN
YCSNxHztqkJqlsdcGLXFxNMTE/2k3ODOiL46f59Phi+Xyg44tzFjb/hcG8q07V46
/7TWNngrvn/8bgpM5Qqi9sx0LKa1j1QOVvZgzdBwvjP4415QryDVteFOX4XpgN0o
ba69lmZXkTO8gvZxpY6RtPrBhjUYrpGgajSF5GEFZc4JYeWxjD2JweGM12YQ3IPc
vmtz82+nzsu8FcAF6bny0hBaW7FJm9HtXbIzfwxQen5a5O/8KqFQUiNGHlsgfS2V
lKYWNAn+8x7LpzRI6TnopfgYIW7+3ur3I15rofWLXnyHNxlSA9288St40Yj/5fXA
OWwbnXZDMB41M7t0hobBhyhI715ksmf5uxIgQoASw+HIkPImMXCdjBlb+H01dQ8P
J45yZlApnuJ+4H6BeiPVd276F6pJbRPAm5LJ3zAzuj0FEUeJRWqnG0AfwnKEe10P
owOGkDqmNwRyhaBP73Wz5FvbIfArwuyrXSvSxtLckZG59+3p1zVi/ChzX4L5rs1W
s+hTUuTWEnAUlRp/TPaB8KTZaKm/7ko5+KklelwbCkmeblgBL4v4y8rD6GjZNbha
SNt3JrT+FNGe5KHm9+ZsZ4oJmIVyDL+HnWt3vjiZT4TB1INeIHjhVwOcrcttSe73
J0mR9AhVNFB01hy7IsaPKAfzI4avzIfoI+IN30elHWgrR6/Gk/ZbOESFUEqSCS/k
g3QYDKpa4Ja5pjAsFEsRZDq8w5/x1uPg37CFnxs4j5YGjN8dDB0FP3wKQhaB9r3w
xWMR67YUaKl96McTLKeAbgAW0xIldOR0QN+17AcLk46EvXdM0Tht2HZzJdkYYiuB
40JKdzlZ2rB4aK/tedQzpalTZO5Pi5ySxbQbGepR6N8P0r1wdHvlm1YXpsdi7gzS
0xSb0mwT6vPQNZkIANL1gbrToxLxYDatqzNlfdJhBoQTRMsEzFwajwLABvduh1K3
TPois2QqxY9J2qO3f5D0ze2gRodOovzioUA6rPXrL3uJfE9bGEK+1N9/x2kFNNgq
Pr06+OeJh0S7GuBLCi7ddLEzZeupnetjFC+ZDbZhFVDLCSGEVYnbe1uoh/UHKSUI
1KNqh3DluHbvjpocsl47dXSyexouPtpcrXSe3yiIHo4LhkWEmopOHDl93rAwX6q0
4Kesc4xKd4AdTKZXRaBOaeP7sE1NdkM3JMJw4tfBpQ8p3EZ3ebL8nMgePC6G9Qpw
LE7PkTz+fKHRZPnHHAaYPHvRVNxBWeMiYj4s9WeXgKYRsVnXGtm0qYuTMVUoomYw
g6ByPspiB4ObRZPyYs376HlwWZ5C29ZKwZDvwIKe4zNxLpOSciRfLCiNKuH2WZnt
5mj/0zRToEfatWwGZ6oX1nvEs+rwTt+Nm6+frm6uW3k14P9K6wyKEors08oHomT0
9O6/YHtJmvDRsM71h2q1Zy3GTJUa7s0JZY9avnDEyi6+iO9ee7a2UGwwft+i1uC8
1XG1IHS5OoMsu2TnF2T26Pw6NPDgbVHLmKPXbIU2v0poJs7PYvyzU9f1wrEtk2PJ
A79Qiiu2JNlTo+iwOf9nSYn+yg1Qq6JN9CC/XP6Cg1LYUpDIF4aCGfzx0khkJAD1
vCZG3tHwIlv8dMXxOnYEKRrqhgT0lk+TPTXh0/L0k/e35keSQTzawHTIKwFXE/rx
XWHwJSQB36jLXNfKOgmIg12VWKb3vwie/G6k12fTWXN69id+etAaD8QGZgaDHH9W
C7J2TTjNLWoa25u/qMC4nJIB7ejZRKsNCTcjOKhtteFO49Tmfs7l3w2PUokl4nWa
TbSRGX7DAEOs38VoGNZTcPUiG3wXnugy08GJOlcnwYbXiC9sRZG/chhK2D/V2Vue
i+a3vEHqEHbRU6FXjWG7s0MtjfIjdBQJO0XbtoUSDxOkKTJmfxHsANdcCvbfG6J1
+RmoBWtPRR+CFiJxcvZ8nfrkWomUSjo0X4g389qVXJ3K2ugZsRUFOvg3VZfhYubu
Gu4LPvKhPuTysveM4vYTAn+fSxgzPySt74f5AXujnmesUnJT98gxXM54y9XPsrWZ
TwKunYXmBrOrbLz9mDowXXtIa6OQ5PENO2cRSYCFeVNk6ekf8tm7FG4oqv9gR0I9
R7/ft2BADsViDkBqpeIvbjisFhk5LxVIzqR88Knww2Zi27KrTgu0/v8ZtWwQ/1tr
3vPbmfgP0m2vJNyLibMUVl9J1flnWB92keo0HUlgVd/Bf7ID1NUEXfHAxI8naq8S
SGQ0Ndnyaq1OQy0275hbm1cnqhnfr8Hn8O1ccmRGdkiTOLlECrzKaRvMPg6zgJtk
sqWrCsLH31pTEaa77uoBdUtcVdXp6Tz57RV6hd+QsS/OKXFp4Gj/JLXSyCJK59eu
4bvfNGDJyNOD2LCJYkArHCirzGe11QqfMQiHWibcb21rv4Bc7MUJWVaODIxPi4mu
B19rYHBCQ3f4yNjCnyMNwgttN08DBdxKJRLMSprlLGcAZCoVDmjyiyFGuCA6C6lu
kKoSZ1XsQXqikboAEMTlH9nHkWwwUL3Ni9V0z91XJwRf4KWwxNyqrfmbkIU0io8D
yQGJZyXS4IYqXv+iY/sojg93YJOcRTwueaRTNAztBlxIolwzlFRSniGRqTsShJtV
PIZspj85nYuJ5NdIjbRRaKCXM9nLL4+0B4CkeeG9/E/+lgDS/6bhtH63Gef5lOto
KDWq/oLnkPNLh6FwyQJKKnaM4DuYiToHVssLkE85QQfY/M1zluYYH5POD2uKv+9S
qFLBLFg8xHoBrHp0NMGn6Zo/zEGo4slv79wB4N9uSyMWIQfmWh55Cvm3UzBAdLx2
3mNGAPZzNhfPsEzd1XehAOLkDF5E8JV1r2D2rn6PsaD2uVt84etPglpj/tDvdxzz
FHlk/Wodn/MzNPzNvqO1bno63yMr/j6WMv4nduiqsx1GB/NXdI3Ftowb9SEbj9Wl
6/0PPKq8LnXE4c5hVXFs0gmA37DxVn846pHYv74dRbuyKKtEqv0OVOT0eAzd7iE9
QZbx7hpMF3GFj5uPF/ClIoe0ptxdBbRrRPdYNBenrmsRfonkalo9Iasu+lle1TxZ
J3AxZbxfyott/C3MIi+16VKXLnD0Iuye75KB13FFzUGSo0ewN4zyOHbFoprJh4To
eWHl88O/SQSGijPhkZTurZbPNnrCGcKBt9q9hod2hOXyHcxBmMOnPGJ5V7YZI70U
tBLybDzxu4HRCs+gz6RYIO3yZPLb3CpnRvbpuIe3aB0BlhoPQpvOqJBl+fNVVVQP
pgbYuIFnj9Y+Fh4gm0diEcHjpyJYSvl39otdAisdb5qnnIyiRN4kpE2mwVbkyCHg
q5yCRxYcNZSiu1XWBJzz/urs/kjFKzobVtFq7gkSEx/ifGM5Px6oBtnpAYHZA3Z9
AmrETg7cv14a6pOskms4Z83nzMaCBuRuWR4YOB7HOxwjWXIBeJKRl92i7PHc3zzd
j8p9hDkf5KI/RuUhQIe0fW5zePkDZbVXn8mTL1tDAcaahfI4kAGXuzhDCeBcgAYm
yidxT+8dXNLZk6xl5tI6Kc7bwda/HlYqNKmuYxiexaZZltWarCibOvb0q8i709hq
M8dLogO9/IGChaBfnge6hOAbt9F05l9bdscFUvpqPMlu6d2Qs4PXBOYaJvDl5bjA
JBJkEIm2iOslu7EBbdaIMTsd6YN6dnrIISaUlmjlDBlnVXDvVvuGVyCvPDHWfI2/
vh2eNcL5ahPwkWDLVODd5RxF03Oq3EoV961I4wWpXr0h4jJJ2MSp4EBWXvx6TqY2
qE3HXfTkJvj4zNv51SHTozKZenmtz/wCYzgNZKqa2hSjlCH3+1T5CZM1SFbGdn6q
o0itI4E1hSBFsYiQj2TZ0sCufmS8NL060KaRF8V87oHRlWIPo5cdvywjUk5+5EAr
ukqbK+PW6Y6lHNO5pDovCI59my30FiFYaKDxayrZ3Dtxix0WR544HQ+CVZATh5+P
xtdem9g0Hto2+dYZrX4YR8iYEzJHOfIH+05mngB+30malBnkneIxqXZxtPxJz2Ac
FmboavDwzloakJ2az8s9/+voZaH2WZOjGBff2cepKUkRie18I6AM9mPe331S3qb/
5WkoqzGipE3VA9otmEavn0j+tTa21lf6DGSJb9i+CMb5U8CtV6kNDmak938oJA8y
CUGrffGfzH+56wlFwsubgJW0kyE2g8W+lb4EQ4Fk12eI3/EpksQOCWQPCDs0OX7d
n0ztL3PDht47vGp3QvmVn3IQu7jVO6VaBaK6+xVUIUdkXYnNOu++GjHP1brxBgRH
VXUDPgsljd1UI2Zh8K9+a3dIpNgKXhxrwt4MYk6Elx0Jo0dS5vb4SOIHNB1oLryZ
LdRvpoQ9hBAoUMiCTVvYfTUSs5amTKlABFCMbEHuHgm1DlATcRlMJ/sIBetsYuN4
3KT3CzFvmo9Iby/3fYlVdagwWdW0wwVRo2HGlLSBYkbqT4LguRbAySRHOx5Ay9Fy
NPz7ERqUIMQgvmO8BmcHmhX1SwszQldtIsIV8lD4AZ3KMLLpxxgCN/kc9jWesU57
lVCM3GYm0/u9YE7tulhD9nRwp93LsCPv8HcwgqxE/wQjicLrRJo+8SjvPfAqY4Dg
x9OGO9tvnx8SCrXplCo3el09LXo9nlQzQhOpGJMyDHiEgbCUXz3aR3ZCOb76i1Hs
JwvP50SCRdQG2OMCGBPI4/E1725xwZD2vLuPp/ZRYYHlcAzekNmn2Gp7iHoTWBoK
ChH3ks90WGCkg2p3t0MFBTVu75/pmrn6VmJiQ/kzkKmz95SMjEf5YDNIae284cny
BwR0dnDwMjDjgflIdy/esZSmHPqtBIlJJDPNH4Bk2wRWQnVKhyy/x3D4DNAFJJKI
SX0HPAwCbko7L7UpuvjEmuXcb+lUuiEXy+bYWNmq+YJxxlOsFprTlZkEABRH8bBL
pnH9gA7l/uV974OX7ZJWqNWTVXzMPVP9JXau3dqnK5XJP0N4umY9ImXFJj7NFQf+
NC3dPNxep8484Q2v5nOQ4fCd1NVneI5PiyWA7ZCfmht+VGwwGRQP7BYpnRp9syP3
cIkEryU3oFZtYCVz77DOIZWzcNqahN7f1Z8cck+X47Mf4DZXPh0BpMKirFHhYqar
QnYr7Bqw7jWjIy0jgkWabeG7m1jUyzZ/amt+/7Yg33c4BR8M2EdyQCVneKcqcSNp
INHH1t0bbt3c5NbCRRAeZ5+Am1/ALjGJ+nOtSQEzt4Cbr4rgwXg2DuaW1WyJnSue
sUrOHD1dc0u9haRX1hLzuVmDHyN57VkFuENVogq0s7cKpS6lnyGAKhru1gvtrb1Y
NfM1aR7lgIwYRg5K8oHAJox4iLhZho2qUoF2j570fERLBNyczTnSpALq65iFbYey
7KiJ0QGcFApBLZojQEvU4TUs6AejaQPTsEGnE/qyLAxQ1844bbq8ajX5HkFosYOz
vP/aTsKAzzLXck/enZ7I6qK6NQiZ4YXUW2rTpjZc+asUj7S3w5eTc0f5wWSIGXZq
m49ihdmkGEUZIwRG8tTe/aar4sGiE5EeyhJ4ZcqyFoea60QMFgDEcWoCRRlXykej
wN1+No99VLAHeyO3vVga/96ogbeSsl8TRtnPtXq2sZ96PynPjiNxiX1JNdgwqrKj
S2SuGQA+lJ5pRrrMwYQpi84xxPwETXnaRhPfhIv+/OsGR0RfbVn8JXr9swwZcbLf
+hmSfL4VW0Dduv6ziwmkGwiZeN3usIIGmAiQJwnirhvukk+F1exL0KGMt3Bzssu/
MOclRIrSnnXQp2bPMA9x1SNAa+8P5INo2dPMpB+0fGts6AsxwqNu5K5BlGZtRE81
cDAg1jrhe5Ghv84aQ9C5bw18ToZbzrBW2qBTEAj/ghlHvTMTf472jgHi+T81sMkN
v/Iy+9yc2wxLj9Pxcb5Nd19xdupZrYYLqvw10Qmbnix+19e2FHxPDqxbi3H0qi7l
Whqbniox7KpOFyUWPjh89wOvSYwyi00uhvWFrf+MOAfi/eEqaX/NF5+JnHIZo/mW
/Ue2frD4tn8IvWljK+oxAM19gEPHb7atAzdIx5iIBN35C4i4oulamXil3skptXs+
KwDpiOPP9Vj4HvTDth5UJijkJ2RY6/M0fJUoF18qXS0rRoW2h6F0oLxGSZsVBcio
FpW2tXcqIvMrKWoe/4aZB//6UGnb4rcZ1YN8Rtbf/odvhK/mwDdIZwiT76G8/gUq
VMG+OK3GFXc3O/kS1Hh0OpdD/qMO973ds4Cx6Iv+3S1pawq2dLQcehuGRmFIt6II
yFOYse65t+AWSHqoCoLolcz8siPjDcZYkHit7ntryXlvrWAF5sJZP+j5Y6jtMwEb
hBfYR421P0qdanqQYdX8MQqqtoDM4OomeUtg8MaYlQ0j47HyOoMkM4pZDG+hJyVB
SBw5R7oi6bmIfJGuBN1i7ZGyHsKarRfkTwIKTKSEk6WwDILr9otVvY1xVvcj3eTM
njR1kRWWweYL8XSOaIowLNz2b538iyroK7qima9ytse8y8iZBJDAw0QAPxv+5HER
AM2uaA27700o59Fk5WgKv+PjGJT/z9m6UTzsqSJTBvj85tkfMtAAGKrtZC11lJz6
YL6l6qK+WzLe8dVLfqPnhwXZ9S44zH78TvQ9Dh3cIbfYxvknhAGJo6/RwaB8i9/X
w7GQ6HAjRzAXb0bMXKaOtyCI0TQW89c5x2c2OiKo3Adk+zbNQOJFzmz4CnINlkz4
M/wzgBV/QpQHUkgG07qIKkTLdSB4JFeukklIjfcj6ZyGKadAnLWb8eHo+91gq4z6
a1qzqtuCat+/KtnOjPRGRtJSi+VeTjYAfYja5YEP9ruFfHmFktxJZn0cLdcZ/lGU
INNUEHEKStL0m+I2Ds6D7tfIPIX++wBYHcpSBhC6KAbJSnYHhfm82gqJnIrdfhNG
yxnSA4GghlGln7zi3QiyByxhs6OZY/JcWaUFY0HG4SL8/Kq3v/Fop10nm/AdCMMo
v4zR1xThfODan8EhYZBGeByEfnSTc/X9JhGEWDtFABfAKpBrRKTnYMUgG5e7l0UD
eCa1MInqK79NBsD5FVcTFynVmyaCRsggDnKqJxmqxGBiz8K0IVqH0+kyqt4MQ2ta
VpyCctJdX1C3Pwb2rHjpM/hgsvHauAgijg4vHcoOAPkHLjC94y5MlA4J9Xd49Unv
l+T5eRSUL9NRLO0sGqg8/vi3vqBmC4p7uGk7Z/CqaHBqyBeWw0vF3PEf9HAS661Q
4qS7Hpb35gsta/J/caap4quG9rvGDIxB+9Lo1j0T59Fcd7dFZGvNggX1p0h8bim+
d2a04pi9RFArBqCHBwQ8uc+BiEQwouHRQVU+JBquwtIhzh59/67qjeeKdIFdeETV
Y7Wr9hGMiFY+TH2/kOXWHIqOTx94e9QqGW/av6x/89CYR87eAfL4LiVXnFs92oxf
9jGDPQ2IlwBD0hBVe/FGptC22E/oHVot6QA8jQMHh5Bo5F+boSdwKKvtXEc+0PVj
1Gc9T7Sw73dKwAcm72x8Kz8TLKrf2mAJ3ON0vPwkuwmw48RX3qGFwi7hezR3sqZX
Al38P+lRlB3CZSADCQLzj9RbO6GiXGp7UDTQZAFtNEDkrNuqZcSDB/xuRvlp1Myj
lJTqE6z4h/H8dJCYBzv89PTTVK2wIZ+fqDm2uDwirFS55Vtb0gEsT8akojNueETm
aYg/tTDWfrvLNOFiJi4sW6Pxax9RyssfjD0zD064XS1dgr9HPsZMKBwYWNEQcsdB
+briwHbii3YFCXykFuJ/8Yr0FMNvCNO2u2weOQoS6+dqatT1l/v4soVFxDE5HvvR
O76QfMb26/QhbYzGNI11zlkPpQp3Tw8TciGNTp9EdhJVQLEpCBAm89nwCIGvdaQJ
UY0+m/DsJ6p4Qjlshc034iqPPMSuUAGV7aIEAWPGCZXJesXk8edFsQ2g2PB30s+T
TALCB+XPs/p+wKO/Dii59RBWYZN6fMYfHJFTOTg+vKHzy0sB5oqLRz6E5YcHR1Dt
Z9SlmQJYAPB5j1P4xPlymeZBAzp3lEC6lVyXHQV6MLEBL2FYuw7o3d1JT1dDP1fA
87fXjGQLHR+GETU/UDitJKPhHm4xHI/v8rwo0zC/naaI5UeAx6OSSjw+s5CHO5o3
b/oM0SXao6fsEG74SCxo9kQuI5HOIAIcL3BB3CJMw9AbZof09ThPKhdJMERYw9gA
sJze/L8RcRPw9B1lQY7etCQc9gdIgdeU2StaluUDmC+AdVwOEa1B8w5xJhQ7c1Rx
h2eyX768RrVJpxCN5xJjdYE8CQ0dIBpjg36CHoHKUk3iRkqwpkKNk/KqXxfLZOkB
/YafXWSSdjlffH76gvxERNjP46FdfWGAoDuvdIR1JaOtyOpYYVkmvIMJ6eEPUexF
SyNXkx+wWJYN5HQxKk59/WAN6oneEtAi23Vppx2Uh1ZXu6nSAtzGc9XuYX7dCxpi
bNd24YP0fhYA6Gr7bxWe38TpNHUgmjzBs5Kq+H/4QCi/K2FdxF6u2u9km7MlehGs
MTpBawsAoFNZS0ZoCqDAtpqSs2aMiAMh2OAhDsyFjpFkbN5C9i8fQzT9DKI/Z4T5
6GzZFMUv+QvrDMDYCftd8lfjlhQPOvSUEWsvXfIHG/DstuU5NHQHUwR7yZotpaA9
uMrsRg9hwgGA97My809kOIxz/dAeRPT5KRQwyy+CP+oNPw2hbsfhIAH/C+ti3vE5
Yx1r5KBT5KUxDPp9MkdBzHK3kMydA4J7CA2eTA1tDiT7B9pu+cNHlg7ymTavX/J4
ObpsuyYwzYKuDcbQFyuR2mQpypHXPJ6l9MrAefcJf82biMEBhFw8r0iPpEosQ2ID
1NQpqBjZz7cvAXqJbFDIf8hSyAm9QfB+uyJu8zLKQh4VbqDBB5LKkkEhUjRcqEUF
ZWuoolIdK2WzZK7Vvlk52A9i0O+fuNKXsDa/VGZdL+5I0WDWAk/PjsdTUYy/lsOH
84cgR9VUmw6+ifG12seagSiTQbhb/fJinzwhz5ML7924KAA2/47Th9chcVkZ44x/
pWXCPgskn/UVJaFEKOs3WlqrJvD2sOO3R5PF1sKziMTsFXcEp4qpHUHMRhFQGglg
VSjKjsH6Hhnj/slL95b+mMGb1oSPI+MlYyCNSJRLTmja3/yCVkD1dhcjdn/Gg/V1
cUJ8mPLNzyVRLyR4UY6xgWzYjcUhM7xIo2whRUUW2S+GW6Ih5YG/IZE/AmEMsG4A
JtbPvSsXCHp465cKF13NMn7AA2Dn/4+1X9q8P7AVN4g4aY0y+bfqdeGay2KYUB3i
q6tKPv/hEvZrls5tYBCQbONSzHLm0nOqmWYj7gIoT5k9mqKLTq9zBDSef8thjqAd
3miUnvVD2gkQhv3g8dYCwx/1l+YZ28XDef51hYxYxtXESJbA3lubDpcEXo0IoqwY
HAO/QZPvOZTG8y5bzO2YnlsQaQ/7qmUSSl5bFpLXx32cpTJK8RwW/SQJjDdRUUu7
12QlGNsliuhYICh6XYqR/tEi8/qc6OFlMJH/4oKweJuzsFWBg7gM/aes8bUM8DZQ
ahG7VpEWrtlqNSeqtNaSB7ThSvHgMKcR9gmbzfhHAcO5prSC6YBMfCpUYfj+ACZ6
nIJwZgFwov2yOIK0kUpRQKAesC1dZ3PzbbwlsM1HF6kTWSdMIE7n6yPg31RRg0NI
HFi06kqHqQmcA+1xPHi2X2F5YTNg8WFVZWHyr/mlNhpIDtOtEaGgtOrTPe1IZvUr
fG8t9FSkuynP7+WLLXqGcFMeWtTKm8uVgdSDa2ZF9CUO/xqwaLPcqFxrHVhO9Gcw
l552VxvR1hJUATLzIOWJldTecprwrBGRA3rDlTk/vztWqe/T5K373SpOoi5w/vBK
b4s0WLM5O2WPgibHrWhtod8NJBIjQJHj65cryzrhAm1xH2wyeV1c7Mylo+Bf9o0+
t44Pq5G9mD9xbYvFGcs1RWlHgAQ/bKgRdTi69ZmF9NA98lbEl5C4Qp4eJP42ywOx
IbXU11jXREvQzdEH10fEXhM7wtvxtOSF6qMdIlUl04SKLCp0ISnPZsr3X2sjb5WL
QAJj1JU8ryd9iRdABZKhE0B1A1xvD+vjvTtVJB/MZaufvVVogLSBuUnGK0x8H/wd
arkd6ie5EEoJCN0NLxK1oaS/sDyGYO/Z6ULZUznHw2nKjTO+5yO8KpgStXJgJYYN
mxwVHMZq0YYwXL2smO1+wvBocGoARahXP4G67WlwjRgdquUsF2nLw3+PfBOHE722
9z1BBJbXKjx5Faz4RqDfVa0YAubCft4CVQe+5l5Hfp1bJa7o3cenF+493ppeIbON
bwGoSp3GZSTH+L4JVrVC7+gQMIlomu5ELGy42yLTRKKfCtXvIfa6NC/PYaKQIbiq
mULweR3pNOEMTWicZnSFkW/3atRWPl0wdNxAyUbKjQj89wJ3uyp3oiAIVU7aFe3O
SF8i3siaa7aYNBaKaZPqkms1MR4W9AUUNjSgHluC3sU0IpI+FzHm2hx4ribAi3s4
0NSMCRlcOAvesEjizODToWUMTP9l+F8WEgAJRZgyAYn7xWXDO0HkzFsCTtmbkLgf
vpo5F+DrA52KW/HVXZxYHJDTlgknNZ9oebISWuxGZexL1RvzHxQzhz1cSzo5uPA6
PaizISyL7yFN9/dXzdUF66UvULo9kWjZUPQjQAP1pIbrSc0fsHLocWqBstQEymRF
NcjfhZBv6M7TCG3lrf1uZ6sQqN+7RqN+n7P3GkMFtGnDoqXIGuktiur++xmyK44q
WlCbmuaHr4DraZ8tkD1gH61pKDjR4TsG8l9zpNwRUvTOpzBMiW78SwKryL2+0s9M
cH8WqzBi3MTj9l3QYW6uVfOcd3GwAb2yUFsoNuIcPamUnk1ms7GZff3Ib1/I55ZT
+DAVnNbaw5JOQ0B18X+srPaKoP7KtscHzmjc1kLw4IAH+mkT3DkT3wMQUfTpypIi
8ypYznJkKaTkEqc7vinGM5+DH3WwLMUkjiKqXiTs2tK20BWAHL8XHs9NB9cBj2xD
mlpA6Vu48H6OHQiZUb21XbEv4NwfxOeDhYeHx1cDa+rLxm+tD+auQkM0gxCLAnR0
5ZgKDpB1RDd/cdzzCYWyWI5FK4QLLhb9/jcR3o2MOB0rzdrOZCS2A/4ccw9zWUQ4
QWp4IWONIyRZyD0sY/bcLAbSjTBObyXWeagLwng2GCkrNcrObUFVper1mGyDShpv
ywMvvV8Qg8pQPQARHZ/BtKEmpvGIP7xkuWi+ftvjrVIw9Go7IB3qgRRMddH68E36
pPtXWQLkTdDmNamJki82xynDoVcaJGpp+mhadJqJ5hcBJWUVwk8jAN9CM4z55V1V
kwUTGGYtwmnU1CVoFIis4aylKNwjuXtc3FUZHwj/P/y4bg1s9zjTwhAJrS8258pG
1RVhdqk5OD5K1fMD1LzfM8Y+U8EkPh7HzYCH3EmQ/JcZEZOc9W8mDbHkVedozKh8
t5Q81kq5adcu6OPLlTylcugR77t2dOPqzsGePJfNAjek8iZOPVqJ7JTWiMAbmABM
L/mZq5aHSURpJT8vhOUgDti+2gB7KrAVGdV5+xEG3axsu2Qiy6bFXaTOGxTeKm6+
nj6Mj+upzwX0uyfxLHrXJYZxp8b5yPgJLtj5in8HqK5Q8nbeA+7zSFx5iKkoQ+JM
1cY2uqVxi+O5zcgIhIxH7JfVZ581/7aBKU5U130FXM8iac0AC4v2LqLa3yXMuAyx
mK2heLO9lcbqE6livHVU+gzGlOZUoge+/rzv4v+R3u2M3IbDVEeeQWxcJt8Ql425
G8OWZhJV/dGN5H2Vrgh6QN2Ugx5I0p4X45MvyOrKh/+UXTVPbK0rIZf/rOq/pLer
Rp/CQ8mpsI/7cQ2JEwhS0qfkDcm9wC9ApUB2KIZU30u4dP+W8EoTwJobBNXXPuGJ
wJRQYpiszdIcvv0IT55L6NNp56P0AKsITmwg+d+gtS87A/TxcENJxHEaCedel8vf
/5CZSf62XjyDIkNuSU6viyCAqCHdL2HqfjVmlXz+GV+x/YlmYKk7kroh+zwDFkDU
cMnAtNrJBRR/wOU1jqYO5dEAbkfAdTP6RZViQQL6V46dcANmyfQwNv9wFA61tZui
hR8ttZK/2ExoMNzSc+6AMuMw0BRNRPQvAla9/LK6WkfETDIm6f1ZwDKB2ezZ6FS3
3dj2lV+4uDWhzGgHYXZVL32BYJtvVk6WO0S3ThLEw5AwmbPoidyLNU/PXaJ48FvB
mQ2qwTN/AedMNqTsAMyRy6k6ScnstorxT0M4i93RG5IKI94vHS94Fwx8W/5u5sj2
vWgwkYAUIFl5Bty4DMBpIb2kAHyNFVozSq4qfBpk+YCna3slm4G0ZoNIgLkYC1L+
uwB9LceA6uHSWdRmIRO/oRn4eOZZcHdOMMttgfPRqjdK816v3BsQTd0tobPvm5vo
y51EZqVUY94gnc5erX8fTpo36j25yND++MRPs3loZl33sGcHLGBCmPTEV40070HJ
TOQopCWz7kWnwIQD6LmdeILE9PWAZG2S+yi7zigGfEwtlVPusRiOtx+E1bqfINbC
4mL36g/GMfr/VR694wSHXCkcrCClb/K2usjgfnAu2cLFqdaZ5jKoLRNNCPnpK5bE
8vO98LlmHZpTDJZjzeYkZohC0++2rNwnk7FMtde4LzG1ir+fSPw19L0Z68WuUUZA
0ZCJs2yxYtza9foI+0BkJ6CRogctIL4fwUVVXwX8du9EwGoMmylPZIE6Oja30to+
DSnHcHFv6p5ZXTr1l1/vZymC9jqpcZdyhmV63xxxKFxdgxlWVTDnXUVf6BOwpVOB
4O9uwEsj3qrUB2h+5G5WFTO0vZa5g+lD9wd0rdbxeSZ/9H7d4iu2w36HFgqywDQh
32efeDdIpIhAeQ5KWpQUpT+n/RNL0uXhCOL8bX96oKgCRtBCCklunao66dbHeMuR
rsslet0WkYvuWpcqO0zVYNhyls8ccFlRRPylRcH+HaapuxYT5ogRayGlQhRP7Fck
VYYAuzZgPHaSVtBnQjs7/MXz5oWA5ZqHwHuKvxXPL+HouAvIAEE6iTqGYL8ZT6iW
OTJ+jWvLqcCeow67z9gpLP7JIG3/DANoIBvlOfN3AurB/nPkqlQAuDOgw7BTX6l6
Jg3CPsUZ3wjTo/3K/98SGvNYR0qM1QR8F3VwHauuvGEwepwlvAVZj4KTMA8msL+k
JopCvhZqQ3WcsYNwa/LSnvREralXP4PCKB9kyC4vGZJmZOUujF+iZU/t4nPNyVCM
/LDR25Gbpoo23QG3gDZT5+p4v/yO8WCXi8iN0QU33k55bN3H+YPZqYHFt8nKdcDt
NrBquvnYQcsXa8dV3t63Mbe3b2Jsakg3TYT5oGReMd5Bz1VfQDyUgNG3hExA1RbB
+uC9HzIbDX+A0m59HnNkZvUUjs9q5q+ZmGYXoLIFOzZbU3wNK9RBsAs7/oY/FzRW
AsDoTt/xvW68DX4DGMGaByriHKA2YXikrMIUUUhtNNxNb+ZOkEI3gDGVDw3AGkoh
p4Te/KRneLkNzTALXeV1uKs51YvIHLJskdYA+hikgwUTl3upagUgXjUsvXMWNKuM
6eFLIL2mIpvHYrgdsfmjOe5ojulvehh16id3J3MgNgDWftoYLG9KaEWULUcm3QDv
BBI/rEvQHIYW0FHdddTiihB9KnAoyiwQSB4FXsfqSqrubD6lPakY/MldBsckzb/E
2Jej+oIqGa2gdTeHqswObek+iv6ToSCiVmcHw21SrS+Di+joB17R7u50TwVm6Zmk
Xkd3u5oc3/iSSoIvEnWY60YYcrmBYHmhuriPENHMCs5u+To1ay2+e2Aln0NSXjP7
N9bZfnZD1DGpSqX1wfTmBqOAm2pDB2fzeu14us1FTvVzEAk6EKl2lly9jrkBDfwV
mxgCvYKjRaD3r+3NclYjmFU6bhHcE5MNFo+at0CTvbSGROLaveKT9FIRDc7h2GeE
qOrrePdv1MQeMK/WFxxDAnG6LmbmTMHI0F9JDfNIdJy5bGDcQXatO7xtfpvFPdwT
BTpk9Os01h315b9ZAAE6g2ZXjDGk2gcgWlMKuGCWSFbIZf2YjySdPPSEa9G5+YZy
CSN/+STrWJS2DAKYIBUyIRik1wkPyWGPmgL2TfnwXVEzJlzX5mODMQmBnbzysN6L
jP8rzoDTTA4spv9z5vvN7gReBj6emCqTflC2jcspO/9e3e2M+qMtkTvK31CQoEc4
n75TEdPDInJB10vnTCkJKwlnUDWDmq6cslGI3AUgTG2CwlaSvPC6I7w+hFAwGP+1
AOo6gpgHZbjl/tTOxMSxx/qaQX8yNSxoyc658oh2DQMx0+Txk99RGoif4D2BPO6I
yCslctG+Ll21jZEBjCR3r8r0Gu0oVv+kHfqjTaeo4HWLOrOLtWfemjAtvOvBsoNZ
yjpIdlpau6IzLyPKBPmR4Z4Ec9+dyEo1/pQZqJ2ZVd09Fa4hDyO+gezibR3zv1jk
7pCx03bG2qdT6id2nXmQfR/Eb0r56RGUEQoZON5pZZ3I+zOscxA7XNmmY68QXd3/
7fe89WbAPs5m46MtVMRGnD/6D3AZVptohabqX76RaYwF42s1iX5cgNn2ElScXH3z
BwcnkXTAL2Moyhcfx7uH/40W/TrUz/jJoAnpLixzPE5VL01ojXaBxOn4ShW8mZPy
sQgRSURSXCYq3L02fe4fSeFGYBKJOO0E2EP1QdWxNv+VT1yjCfZHDFcYSerFKt1J
GYD8SBtxXf+6Ud8IU6REuZCasL+uJ8L1T4IHwpmP+QOHwmRppq9EtuMSKR5YwEHh
Ku8IJ8Y0nTYFRR8HfLdJPLmL0DCfKpzjaFf3Kjr5G9nPsdhSAIVSs5zzmzNCXxcy
X9fgDrbI4/U93nn4EzQYVNvMauWiLWCpcqFQbVYWtVlV2JenXcv0wsSAwho6ACac
yg5u4ebcJi5lcZRYkaVRxvzjhm+5++KCu1o+i1JjI4ds8Ki8NHFee5alk8O/hJaj
EfEJuvc4AOd+xhppsxWk4cf3MjDUJU9XvMVrmw3dXr/9+b2+E08hhOZnF7h/pUmk
sB0hH5g/bTbpZbVHFUyaMiCtvRehmK9xhJ3cMX7exA3ZG3QMXBSQHdAh7lNg/4Rw
bNIxO7Wa6067wZGkS3rsPp8z3PRk2wLhjV+95Zew4P+CPLPsf7o5bz27dPlVw5Gc
IO/WPKBNKyqQgjFZRcpZESkm+feJX6RM3xP0GH+470OvwgvitJqEF48NsgUcJCtk
gqDhkoRDQ8DoEkgT42vK44qgCoERKQYjwXJcHuv0S5/eRhXjpIrO0yZ1Z+ZNp/Tl
3CQ2lYVMGqyRTUDUy/usIxjOS0BzdsXECRuqyGMD33o4Wa1OFGDS1hH5fOjezLpK
GBXYeF3q5nbhP6CVdSE5xm0ko/54APtVlhpp8oLbupjpfeO4ZF3LvrsibsjgT5uV
to/wrshS4CVLY2k7j+jwIqMlt1BO04ETLcbb2jbUj4gdK/yAgyXL6Aw0t82SKIPp
3WwNXKGpwUQP1mW6iO9tUQP7UZuFRi+X6Pz75Cm2uP+HF8kbfAta/s76ajaPJ4PQ
SIaLUy84zPoWdS4TXlwIgEA2Bi8c6wFT14T7Yfk0P1q7z7t0yigWqQMuWNUNOnpC
7uJGa0oRib2naRSruiGaO/YJdtnXQgltohT54W14swmBxiVf6dVT7tGIFk6XzM7T
iDX8dBqc67U5QObBdFNwnvUeEF9bWuIWT+rfd5epMPO3kTZYzcwEBuxhlj1F+7q9
7HjmDOO1qQXwyJxiJLANzszlzs2swHe2IaEMtEK6Uxuec+2EVwg/AVMFNKc9bijR
iHo2a5bgSLq/aGRwhcCdWl9Wlp96RnP0KkXc3Wf+Q6O8tDDXhX4j6tvYJuhKax4j
zFVJgEb8x+HUCqgPpiHVx093zeASMekn7zrwz2AzzT4W8g3QeUmeUPtxxk5kbLWv
H6oV/bb9vVy5jZmqil1ODrZqJi4lZ9n/ByxyDB/FzWvJuHDhtNzUzsncXlVLKkVz
Ty6C6JsHtTduZFdYkxrUU8UBgxO6Hh0pAeR7iGemYM/Ae0sXscH9amsBiLV1DniM
FTHvI0dNSP7tnvx9IEsPAaTNvYdTbmcsvFQFPoybl7QdudS9kM7wVrGzi7LaMr14
ilc5LvNXpnNYU5g6ohZzyPyej3ZVoo+ObYZLL0+UaL9jMANlBKerKtVXxUrq3h7e
buOGyBZEhEiQGt3njgEIUitnG4B0GFbA2w3FH5eu87ccuBllJt+c+9NbFuZ3tV8n
CmveY2xVY6swVOFOzR8nVOhCpj/cl7yqk21h96gMiMvGrFcCVSYH0h7sLgsLyzm0
zqscAS3Cq12PtYT/6wACUwBEo3GjWA7P6XWCvfJLDin968Lk3sgM5N65NsX1WAWC
TO+EkClWhUTwcgYCR7/U7+mOMcHf6Q9xUOn7a88mozaSql7317rcX/pBTNes4who
h3cBClirRX8wNNNBl0+ombdVRnpzFAbelOcsvMzvXAvkevXS5H9wALoNIibv8x6O
+VF40rAC8VV57cUo4DuTO5ROcIe+c+j2u4sIKjlmiKnUs3yfcUocm5tWQ0t1gmbQ
OvgCoaTlfNxfvlmbT2cKuuZiDrEICkk7ncIaLeJu5Y10b1YLixaCcLMhjEGqJpqi
UdSkQymL8Nl7FlWm/kV84KNVclp2XYXGzF8C4zhrVtihdbysu9JLBbPpJKTU8U15
zKPnDulZ1HoeQjHMdHl3Jtt2XJfXPv829TzDghHnr4PhcKYCyNI8MpgktHhHH3b2
P3L9XIUnkW+IhWkFmAkPDGZ9XilwdSN3/ktYqEQIcEZFSbGFwiBgX3II7eu/yApR
u5uuisV4waTIlMmLRUtnlqKSSqI9l3HscVhRDZMHZsZ7RAa+6RjRfqlL4HFgooFi
UQ/DPEuA2qqykQYzrnEUovSCiQMWu1K6f1NNfp3ScMUiz4sMOLZOksH6JTXoZzZ9
umbvsM8fFde4q+v5+ROXUPvQLBkoLgDaEu8r376guC9h4WjN8XcSXJWysATjLlCA
0a1+vzChMEotbcKkfWeUMEC2M91QR0dSVXnQ6JsI0FXKS+2LVxvuYJzTYMK+99Mh
EUdSIxbsjTPlRjL/N732vyFL3lgQZv2wQuAzdE6d8TnOxxruwusjIjRH1tyilO5Y
THsERGix4/iXdfhQjG8UJrrHlDT+uJcp1rkH9ftAiRiMvOwocU0TPkZv3FiY7mlC
SrpiWu6sfT84D8jU9T90sLgM9AyJ+y2g3mfSPBj+AvAguHIQYmSKspeB8pcDJLSJ
nr2wix2GbG+YQ6Nog7CnH68hZqNRyVz5l44b2Wow6jTrr4TKuxPg4uweZXDbT1sR
24fkNq767ZwdGBFoK+FCmKUy1Q4jnr9QxjB8he0ecYqXWmv/VQT8O4wneM5Ah1BA
sJ5iPDz7qoqv8f8gzKcXlMph16NegphYLguGHGtQnDiC+0/O56BwQa8ua1IkoM9M
DCn8+aPJmLrl0TKCkjOfV/yl2EtwnmXTVaJJ2c3mWUk7c7fRU3X/bsjAgc3QO1dk
1uRQ+nWb8qXKFeRmshBEmFesbDGCVK/rcjc5g2mBZP13UGAkIowI+ovpMrWC6XMk
VwN7IZOy5fHsPR6JJ1hClLCT8OZbNccwqi9HiqqyiLCcJ3ZhAAKkfnHlTa6v+jY7
6ZhbxJ2JE15X21P5+wMlfKgsjSLF8hvTMaLnbaL90Cdl39XOA+F2jVEVJ2+H/i69
cUsq65q+zzZxHRct4Yby/Mh76GYe8X9UAK37BOTqVLHa2xXyWshjx750DPCzDKdw
dStV1ZIssMQNIazRxITaeoF0XgvyGU5/2w6tfGt6ltox9DpALXvZaSTUOwsyDeTk
JFJ5rW1tP11NyfMwjICAG6tY3NbIDiM9oT9czBnkj7cxQcUNgrzajoeKspod91pX
iAB9fsNPAJ5S7wGQQCJFVci6qCgOZosz/6iFI9pZlcyGrpyYEaDuablIksBI8Sco
xoD9aqj8vlsflb5Jt0Ugeylt7MdV5JtTUny8ZxaoiEPcbT/ZXVac9Dim55g5rNN+
5vLDK3jXoEl0qDNylmITSjIqtdN7ejoONriczW0p/EEFISt9At9PIVZSBvreHcJd
1ZeWAY0jOv6E1l8IomsfKUixz2B3wErYUod/oud6s64Uerb4Y9JZYEXV8Ow2S1yU
cZ/G92MwXSpqteD35u3q3hIZARZbuy8ET02np1tARbDqX+7ECYJNqw9SnGQ8Jcqb
PPVpXRppx0lnnVH33kHxRVb7IE8u3ODbNiHIAoKjN8K2/rCdRaspRCL1nw2P2g7l
l3pzx7h5R/tfBc9PGTDZ5Dkv2MISBs4YtY2X5wxlb4hL90mYEaQcECWPeaowCNRK
QrJjFz5zn/43OKcZE9wTUBEeN2xzprlUdy+jW83z+IKeh0TEzbecyCaGaq8QhhZ0
nxbSA0j6I/SLU5sI3VAo9vr+Tpvxcui2JUvBHeP3HeRE8IaSnHmf9sz8ZpI4cnb6
LeZ3ahN2GeVLeEgih+8iwvRS2+2EgwrVrM3eCKrPZ813CbFShAkpD5C2LxuSqgeg
oparZ39TYSoAW0emqcV6PyHqsPU5cdmBAuJ98nfvdn33qNrd+UMguaJTL/ldwcKb
8BFXuDI/RKvNndc+8G6loKQbqNzqj3SHLZSnX6mNBwn9N3INwZ3OVJ09tqaG2x7x
KvJBa7wBbCqabGAoUfc4KKcglQDZAyFlYcLSECZM1VGq0nH3LXNQT2XkpxoGcTAh
NvgFp4bFfN+oCPZf3mo9XSKcpNMiIlK6n0uCRIjG3sT9ARyw7cNHByDqhMqjRlI7
md9EyfSutO5VNUJx0mOes5U4dGGHS8/3MKAgQqhQn4b7TUFr9YRB+DkaOJFdBxz+
RMMkqCc4OipKGvBFClV9twoGRXSCm4uxOpEH97HnJ9iKM8v/8xDdtJNfA205lUVF
AHlKge45ZWt/DgjXrvuiXaKjIZpM+IdcIU07CEVtvuawIsz5LfTbH92yoUdtmcGt
CHfHrPJjG0lb5tED6tjL0I8kqpbY0PXcQiDTxL1HwBi5gMsPhCYZ7BZNuWbPYtov
EgZdbl7YZgYPjaXYIU4wJ+wUWle9lc3K3c8SnBxZ7WDFOWBKV5xG0z+7GYu+zfNk
9X01hJ5jIkbF5/u14H6V4GEIzyfWVQ10YuPrPqoNCFZEwzsW6IfJ61/hpJ0DpL8L
0D3doUuGNWLOSZGZxdvg3ghSfaAo8I5U2rWL+5nYhZw4GKd+MDxEVPyjpmiQps3k
P602qpKJNbTsmvcA8G4hBqdQNI4tjvLMx1Kp4cuMukVV+nmX93SJZ5P296Fcdm/x
siqSEggl1t4bKJTgdD5usdjoQly7q5y/TAt17D7wPjudyqstWFr7xxOqrDu/6JQX
FB70hGxjXPQ1F2j0rckOledQsB32nj15B7M0ER1p/Q7sBZZpB+InyPQaAu8o1cq1
ohrO1kNLJxtJfCM1PhLU92RmKoBe6J3Vik2gVqBUTyvDiN9/eGSLIVXuyAoOTodI
baOBm2aJ3VaSVz+3VGkbMy1IjGKDlhJ/7GsmnPcrwa/XkB5s4ijks/vZwdcvlq/f
ML9wBBqTU/1MGt+Cc5COIIQ7ngACpglthw/7PDg7l6nSOadv40eXCWuntphysXz4
6S75BAEmdMrCRt6G2BUoQ4SrwLBpKxeroxTVJKR5SrkTk2YsmGiQtJ14ZZnnJ9zo
Jau058p6GOmRGDIjVzlWP93VpXn+JIcFim1Gn7E6p0/WW/S0o458s1isfkd30IjV
61BtUs7D2DPEG9ma6khbIDnzDh5+zB3tsFhiKk+Ee0Z0N66hGL4UbWXWSW5kHlAR
9DZHiZQ5swMeMarF9DDOO0T4lVP84FUxCYNRpQ24m0xUjUbMVnxLn7+K/7t5LQxF
BbeJcYTagpe/NGdv/WkPxnBpRPNrERYuc+AzU15WgZ9VUx6NHfylHxpeE8dMjtAm
KBvf1h5r+5iCcsNGo6xwjOb2YqslaX/mKtA1uh42fYhgS+vOteAFDrpCbh7nQysF
4OTRPTkYjCdxvTRDGzm+cgXG/yQ0XHQYjxECtbrK4e2YSnUzZDJ9omGxZNc2B9MP
GITsH0trZqq52w5cH2BWoNLrtKdKrhWOTVFn0fajxkg7aa9rr2XmHAKIQs17B4eN
BPqMJ2jFB+XeAdBRh8T+HfM3e3ZfnLnUnDmYGaIm/V7xhm7330TsbFdU2OHM3FG9
rnlFiCDvdyJMU8dkIUB4HbXuMCWouUH2CfGSh1hJHh7JSNQX+KjP1A85YnTU8SW6
s3JwSdFOlQ8A4JMAX5B924bjEo2wEgeZy9Uj4momGV9ARNbG79qdx7MM26pdTczy
tDKoyAaMtw7ozDOG3aw8cVLUPxW/SMyipLKfbCmdvw9bIJ2XuREB9xy1R068r65t
qCS9oCU6MOnm07LHemzPv6UpdjmDgKXauUeQQ2yUI97z9P9in0rBtVwduFLaDleN
n6evA9ghLUWY8Gv29ywFCw0VIBJKyNUmajqEith5ofCSesw4DQWF6esfV07PSGKF
08F4xjG6l+J9dQhhE1uqLPFViO5tkIem9xQ5Su+rDLJW95WTSbo1qV9ygSiVfNbY
2/IWCc6r5Z70dZGwQIL4zjmwqWslnvi+4nU/xh1NCayVx5k5t7I635qXHsHCLmH/
yUM0ZhcmmMw9eI8fskAPAtKjnxgs4BHyRj5BbAUo/6zvE/O7Pr2EVcYFgSCk9k4s
yW/RvOB2eR81/sRJjxSTBy/xqiXz8M0E1+CD0JGA4pCLeBN7rRXGXUmeD98KowT5
wmNQrC9lhSw5DMqovPTXq/u7yQr5OzD1VUrxXCRGKQVaLcwD/W+mkSDBBoCINkDW
sq5Kg2NdtJjXh7ZKa5LjzqqsmVM96Etz1K8h7CDhmGzhJGxhPv/XaSRVEvrIbY0m
zeIF55Yb8EYwzhFiPDlpVOA/Q7nHIkwCSdKEAH9F0Ig5Wwhwy13v69wQZ1nvsMW1
zazL379zhBY/W7yGZy74yCTVQOGYU1IxJq6uwAYkb3hAfAO8+1bmt3m1L6M+ZUnQ
nX+ebph9MEW9pWKloiX2fLdA6g9gjod4oKnlq4eEFUBaKpLA6JzKenYcKHZJVtQ/
C1lRCPzm85BIgoryaQ5nTFD5jNZjyPKpGWDi8OPnAglybPQqirc6QCsD8Wep8KpE
1avnwkKc8Xco8EMGluPOSQoNlodZQKPnGZfeR6vNSbYmw/RHXNMAhWu/qYyWdBil
vXMypjWS3x8UXQYlShD3OjA8/AajNczt0+QWrLSCj26jnrJjo9cNDym2IwA0XHJL
zWXxfb2WR0ASC66qMYwo4S1pkwmmyP6swROLNEnOSieOny5pM1mVY5bfLR484DSl
qaEXG4CvLOtMCjzTq4/DhTmtDPOEU1Wp2wWT09blyyw/6gmKQPChNgOqdQsafSDT
qPVZlGsG//GbgL3qK6zlIgS90aM1T7ZXRgg4GIYjKj1PsM5rVXXkGIkdSWqgh4sZ
Rzf017ohOgXAcUGRo1UNKgwTM5nJxJMj1YFCZddiaGDUyZtRwE1abaeFQnR3KIaZ
ovBAo0KtAOHxZnj5uRW8pYzXD/zDPu6ge47Hxq1JcV71FuYKCTqG8GciYToUMHOJ
UuRYjARcc6Wur4rIteJoYhb0YIkSIBUJ05ZYqjFSNkhRfb+Ca6KZchNjCs9IMqjV
+mHXbu6Qt7DY10Nn+yps/rXtguBOMeNjccaWxbQKeaiSE2emujJteX+JxVkLwdzX
+g14o1lMFfXHwAjQ4aINVPfrc3n2bYVtg06cyr6pFNQ3SBDo8ukndWwUJO61GOqj
jYerUkmtBzNh8hBhXHZ3LBQu8KtN4UgOgDpu/wthIQoLuFY3cNIxrDh/MyECmTtz
UNV2C/JIsMACbUUGT9qwPn6hTfrIBzvvA5kxvQaIAmOPoynMNJsMh2mjDK+l09/J
n7Yih8GFx3kV5dAg+kn9qvej7q9K2bf3jQXBN0rg/19hpvXYcohOkd5GapJQJyjM
1uD+fmY/dZBFRHkUDehPW4y2oo01uHDaezVLqYJ5WcqETXy8fGk7ytxUEjd2r8Ff
e9qS7X12VAz7D7HDI6GaycYmR8n8Ej7K5LnyfWo0QxS+qOSrEpoVvysw1xQ9Xhtz
uCBDiJfmT4jgxj0lG21XEwX7yjC3o7Xj8Ypy0AbSCBc86edHIbgUmyy5B5qpvb4o
n4vkIxgsL/V/vgq0Q7ryQEkPnPXy1V7pvkfcTZucwY5mkfuWnTk0OdoelxWJ34sx
GAnkAweNIZsdFs9WqQS1Ljop00gudQHKgvz429oQ7ztD6rASYB+Io0BxKJWubIKK
/fm+Y6EXNTDffhJ3XTZppYFB+4xKc5PpmlZ7aRI3lfiz08u6w2CcCNZhaHYp3tBF
SzRo07+uXbhev7GD143Mnh+E2oRybb6lC82vXeaZZ6ZDgO5JWZ9QaHOb4rK5vSPO
46TYoqBMkTU9/g7ssfZwCk6wLvEQnYpTyRlDzBN0F12K9WYHWC5moJIRI+m8zpzU
9py0By5vmVmyWV9P1ryi2NGJxVIiFaVChadZloLxzICDdqIxkrpJAaheRt98uWAb
S68pB+y2vZSRg3ovae0hw0lT1M0BUPCrhpG5pwWdyk/x7+xCXffA95zJMqj0qnZw
OnmlBdThxAGlFlmqTUsJpgZHQz3VeFH+DnoRmM51Go7ebpNonEJ1BQ6oVvdxJzzp
vGvarGyNlu5RzZgtVBlBwdc6fihbryo8WaBqThwuozsQmBVBWksxR3AD0DJ5iNXz
6EK8ytjaUYxZPYCxeQ86mFhSSt79ty1mQtz+k6j0/6kj8USF/9CZNAk7tHmTcehh
zPB98mHN+TcTBWveT5Bi3fUHeHujqMtsV7CvAHs7bZ15+UsUrbYbq7t2LQFxHCQT
gmXKbuNgqH55U9mSlxYXtHKcEtQDR0ylrTIL2XBlZZwQzIYGfsscaGvDHenpaXgv
JyGQ2SEfJh7DoghH4mkvcnkP8ZesIMmFGr7+vOb2A6reEwecXc1XbozfZLS3lRyS
3iADYdc/huV3OL9P00+V3Nnvo8cRDDsHm3m88I0xN/XMN3GXt/YGJGOCT91AChdr
OorHAKSQRXmkGktEGxwh3+42mHwPqvvih2ysp1wJ+n2BrIBGwQeHa1OQZU0VkvhY
SHFjGOux0pmaCOxYOaBGnhLns9GA9NTrvLqvzwI2ob0GgQsh2GSCwAVLXk+nn8hW
FfH/nWY7IYl/zGmot1KB4OLvEdsOi+0DgcTZVhq9b+zShaHj7iJKPUPRkWNEgXnu
5tcbawqB4Shylr9yHgKtZzdfFWTi/zzGZM5/FJCZAqC9AG8olsO9JGX9b97+QidU
xYXLhBGhLb8xJz0auJwmZWUj8A3CsURNyjAH81fH8mD81VVCyZmwWq9E6WBBZcYL
C9gydU11xe8zKY4/AEjUkMs3R00aHcrj+DB+jBj47F49el/tICTYGnKuj69j+3ru
+Vckg8NjtTUMOwOjIgPb7RqWNmLdwPjpOzaZyhzdM0R6PENJR0dTbPsyY5k81WLq
cgwSDQyRg8GbGVwqCenMu/Bt05ML1UdAZihJRIme+Z/r2pKDxeFn/t+v3QPm1dKp
fYkr962JJtyd3D0XMjU0zV/yEbJ2Z+svNkXrtEjdnONSw5DDkvS/eJeZfY8M3FZG
iKaQCxuGiIqC9bqjl/l952rRYRQC48BCVFRMIsQ/W/7K+ru35MR8539CSoD6zNbW
s3Oo0dnoyFhTOp5DCpFk+YpcXn6uuN9sr8AxPNNibSb0MNTd7dREmYAUuC7ztTka
udWnbi5FyWuUwAGPvB1rEvOV7yLqXAbR1g1XH82wlpnoEYmXyXYDTPPlPwJfZPzj
kblqBHArDU0Zt5cOJGgUZ0y1KxJ8rQNr2uoJgcNKuSOahzWutK7p+mnp8e3ZCLKP
Z3CQXPUC0Lg/ztTuZ4NJjRdxHLAubNOtAV2/x6xhNgdyQ8eaJ/gXsGLwnaDd12iC
OwgMfmFtaObvyKFICBe4UXF/8ulnMOjhumA7H4L83cZH7aMaF87J+ixHPjZ/0G22
uCJxCR5z+oOYUOhEvT4Zk0GwWjgh/4r31hPIGfGKjEY3dR564OgZHalQ4ol3LXI/
eJYWCNQ0zI4IIgNaz+5+QxV1s6noEKmZ+fdfIZux7KeA2f9F2naQ6iMMlant2ML7
IKxlxlGEMnaBzjKOLVauSb65I4E3z9udFVdNt0opDkLe9866IBEeTn+WW6b9WgLS
8dOxsb4r6a/dmpCpxD649IDgYNnCx4lBKWroSxzagJkAOKyu49GRzRK4Jj5QQH0a
Wpppi6x1dIBv19pDDtm3xySfrpRWVwPxEFASnnFjbFpJKNzhXf4AVvKpw7HGANHa
kCcRJNhDQdQecxiYkPFTlBDotSel3WYvnttwD8rORgiXPdLJpsadf84jlRvRKtu3
CXyGql7llrVnO6aOmW571tQMdrGOaUfjl1WjEcDEoIelVlyJnCNR7bz4VlvHEHXJ
YDCM2xwOFEm7WYeKxN48sW1tKUNRHVriTfOyxWJF+4GQVUeN1Q1jLk4mTuK2ELfX
xFh5RxiZtXidwJ0b76VYSZkXMZw9pdmgkj/9knK+md23QHlozQYV5bC40mAhSTVD
gxwO65dkHb+44Dl79r2GzZB0xqA3P/uhZ/2znNStfbnE4BT/e7BDhQENSyhljUqc
4EvmrFogli7B6c2d+Qk8DBXqbb3/X6uFbAU3PSDm7Z0f926THZdRgRzlkZiHmJXj
da94FTwOgfhYpFjP0c9WyPjXppOlfrIwQmgLliFO+DcVWQNewIjnyYGKuvdLQlNw
6n/FHdybesxDjJ8/KTv+Hz1HJXLoyUYuljkgidwBRuoDKWMK3eSnJOyrfC5bp20E
orpogN4RBD9yy9DGhksQeAvoRQXMYx4m/FfPtUbODl0imNtcyVGr+I3XePCt/r5c
1YSDZlkZuzAZ4E8b4RjCjmIXgotQOyJLl17jVzhTplzYUyz36aZzTpa8aAIj4GeS
eoMhr0+b7c4Htut4BobJocnYH4cT3rlaXbzNGJZ5H8MOsa8UYTmmHPRV6TYYam0f
NxVPknJE+QlBrULLH3B8+qGBf8bLcskegwpMUUyqWjSjiWtM/Kcn779X2NTL872r
Yyd8L43SI7y4OPxBPu9OoihLrv1eD7nFsBEwGuPCreT/J4lM6tRjnwWrLRU+xkJz
59TknZYjMipuWHRGTH1shEMIO17O5DYoS9QIfKXr2wEGCRhrU9pYERMqWAYeTZ4v
V6RMoAPMWdqCXCicbVdqdugmZAnXnGL8rezzym+Q9ANR7aq0g8Grzot7X2Z6MojY
noIsqi+do7GZyrpY6iD7VTVmpG73Q6KJhd/1IWebvuPTprVVUPElgjf5ezWxcsEv
MeKHHc5XWijixKrQf0WngANkWHMPhSGF2L81/0fyWB75wY5aYBGb0e5mJJllNAEo
L59CHK+UnYy7GLQ22gxSvqFICNlErX3owS7sKXWqVMPiSRZSOqh0hDn1SESO7eQm
d58h9QeDwY2q4wHubGbNeHwMixHQKt+jUuHoZv4YdIf2R5hUyPwUUlaYoPXT/oKA
ztSq/oMbQWuWZlHOGAPIJU+fUKLJ+wBwd18vpkrqvrb2WeyIsCX+JFzLa9Qc1Ksg
oE3o20V1UYhO3f2Gnq3wEwmy+eNeLfYWgvdDFL+GGp64F6xz2AfkCo22qeMpJPcF
hTBVzOyOYXx47pbu+evpKlRTJzvxSfEmwqnT+BgT3fmxdlJBVn/MWverdzAzPV/h
yk4PV1LzpkCNOuT14XgOgboZ+GcEzcpg1XgYv6BNE24MnG2fiLFbwBWmYFTNaeSu
Yryzmjs3hFIhBZOUbGmLb0hF0UHpj/wKJyYvT11sagvwK8eML/9VVG7xXyISPAhu
Hh1H7QDbrp3wxA1gGqoN/jonZstZstdafVUSc0BWxM80b/9Ph86g+QUUBzaK6OOZ
+1BYiUFvS98fe9sEXDXH8v8JGBmon5kE+XOqEQP5G+FVyV3dEwRRzQJNeSi9gYkL
bG8a2Hd+vlWJ4at8otnXsgxG7Ax2J22M3c016ojDKxY4jqvh51/CcJctdrqM3Gr5
0uQ7mw6f9mkidOWkHnChXAXqhxudMOYRne5O6PUcXYOaBBRWSdLLqJXFu5TKAOi6
Vww/eMKqDbrawJhjONZ83TOVyN9F1hriOgsCcVeTKPQZDtoLvOnifprcZTRo5sJ/
fygABw/7rRUdM3PjjzOqFeLCdKiQyZ6sfssgPy4vA6wMYltVhoIr+CZlco16DnGH
eZiB4qd3ullHvoyqI6zW6qpzX2Ct+/Zo98RStITK+eKY770fPvLtD2Twy+E+phph
TsNI52G5k0wqcdBljZxfRd/eK229YNJu0hOt9FDtCn5J9x+DCcBszqbEKM9NcvIp
5k96SWthgQV8gG8io/Aztcom1zZdBxMY0y+A/zRP0Wlee99BcAQO0N6x9wIFDiKW
i+0pLGBNiWYDV1NUEyvcSHPoyAGdFeskaO0ITRDhDOQaHIRbXm2wqzF0Zdt26Jb5
bIgvNVco7EJPYUF8FpykwBY1FAUZrmmR0OnWogCcmGKJjN126B48MYVh1yJHlhAJ
T7RTuYd07nKUFKi+poSJXrz+cB0dmp/dmTetrUwR8HZZ0Bb8+em+oDT7QtbKuSUq
vzMoxzFSaYeiW7Z+bYX8GQZmsB3TgiQhFd4up8rTRxufwsDsFPCDUg1iAo+inRH3
Yc7MFx5wPi34AhbPhyb/Y+W4I/t/1zx35Lwir+8EEqjNB+5qJGilXzNrCjEfHcHU
bdAFLs0uW0JGP76yEGbNCDYTdLt/EnOl5kdwmaYVTg81uz5oIApX3Y0FUCXPB82V
f4POEjRMCpCo0K5r/hQ2nZtVR9vUZ9xY6+T/Uw8bIL369y3CYUQ6lEBxC3uZpevU
Hz1oPAH6WrjV7YB4jsJj7VNxMagPSbcqaJGo25U/BKK+jgpQbCOlNyy0ByURmAiG
3SpkcYLFUnrWZvEnrJEtyebbi5yBBFjrquGecTm1UniIfxrQ+tiBHvthbTOzfkm/
y/QqQTRr1zqgkOspUnt4jm2n+46cLLgJUkWzSRHIOkgY8cxCssL/3+IIZSVqLMOv
eZK0tXqxi5RMRGDmx8Q+bZuoh90TrCypW0s9vYkubpHQG2dq2ttbtY4PY0UIiLiW
ENA02l+N2Br8m0tJY0CP/bpFf/ivyQVd5ZpwH5udL67M89/Xp1VA0+TzKdIx3dCl
YTPtNOuPZyWg5JPEF5mmSEUhixCyuj1RrYve5k7EUzxJNe/9zE5pJc5dQNDP8n/q
sEmdmyURUkLJrARtCU60G1xqIA/IyjjLuca2JQ1jjTpQgb/lQyfCB+f6LL/L4sve
VTcj0uWAZl+HHTfyJCFI5tdctRSEwhrLosyA2FhQ5GVYX9XBQ3KQjVmgcUsYLC9q
xTtVD766ZUMvfvQOG8pPkUv0jgQqSU4g0Tq00vNiOhpRQe1n5riatAKxLvnd0qPa
2gx7wun66e13AFC2fkuCUwctPmtg09D5wvkYXN0b/wn3Ntn+FLlliMoXJ6LAyNjR
Yi4Dgmgva3ftiUxzZaXi4qbZHiUiF0FGR7zPYzir5Hhj14twaoiLErLblmasjt7n
IO+bdZuNBFQ6/RQb7H26VeyHYLuEeRtjqwcEoHAib/5H4YHMMim4zmO+CH5QDNpl
rJOnv+j8zrTCGfdtji53tFu+5bLcxtS9GexNF422hZKVQ/+CYJj/4APqU6fivuNU
okRLTGWOZuD61h+cs/KGRhzcQH90qkDdIUD150ZEw31QT6oM3TPtSBATc8nvg1+X
odw32MhAR2xLkwxbxGG0E7uo4QG5ydhLwnfEuNjSGZXZmY63tjWY/mObVi6mML1j
OUeg5rnOgx7nKvnV5kRyPsOT+cl3LnlqeKndfaoEneWWhPzwplDUXI8P8QigPDPd
RhwlmhfeTggPjK+oFwFyqfb+JYAaKXDGgyF3HLt+GidxNRteyF7K1PKQEpHWmRzK
GP4HWG27eqjF0NA7EsA/h12ff4pDARQHiJ4w6a54laRjm2QCmJv5uHuscYdGNESv
OKyMADyV4mI9P+dMwQ/LxG15aUYcbXTECsH26bReT1qPYa0VQyo1OoQrXNY90kJa
psFnTzK7GWQVXvodMNRx7zcM55UFFJWY/K1V5LpeHfildwH0LKMQ81VfL9UszW0a
ccdy08/qfpk7iC0+IxZnSWNk0i7CzQOejuerceyUafL6BrfPKp5OP++hKDVpVSBu
mSSC7gzNTzZsU/bBxPVk7vKy7U+n5UMvDBRExPqaFj+dotVm2KP/8G+Lyy1Ok4ir
A3c4bOu6I1WbsUXAB4IJ0vgfmAkBy2fNVuKufpoX1/r/n717LjVCJTkanplWTra7
lhzw9Q/6y4M75D0VzOcslqRLLNkd/4vZSa7TESX4bJ/tA9mowC/ADl3TY6JJxGBl
/XLLw0JroqdphgcVrMv3f1PNHZSr+aWqToEBfdie4Kjc8+dNr4X5CL6GdraO+yTt
WindMR7SOA59io7FBwYLJb7mc22kwyg9xpdpj73v1Yh2TxlW6IR3DPOEOzLnHbNK
xStMhtpynzYRBaJTufk15Qa7Sgj5T09KJlBVKpt71f5xTWvrWJgFnw/NlWPf/wpQ
mPsXr56cpngXLfpJpoE/LKDnpRud8j6Vmibpdcmjz/JSWBqTyLV+yxOPwl+m+aER
a/bjFIDih/FZlqqXcXfMwEELOs9ON9YORsXhdwDXnlMHGIRiHKNRNAVagckOEueD
CMGSsszsnDWfKo55Z4LV/WO0Ct6rCyw0krgq3iD7s/lOBuZlisqHXpOAGgYbWa3e
rSFRYNfFFF639/DSoeISvASMZ9dodm2kFBsDJ2uaMpIOWaA/Q9GAr+KjXCra9/Mu
8e85L73CWW0Ut9bPmBx7fEuQtul8KGaf7XZWjJ4lZe24sGDKq2FrSkYUvs/FOaoi
2NjdODbaeE0uxXHjRM5mhhSiVU7twqI5VkJWw/XAdz1rW4JWcuHCsyibuVA9/dMw
DYB+/kubDPb0zm6SNDQGJCIU6zI/aN2gafsTEDL+4AeLvEI4guN6+cO3KKD36pqh
cZNDnjfB/3F9yrlSXPs0NqAi4fAZkjbD5KocVIolGRzDXzThPOwbruL7uX1WfrsT
a36iwEcxxiKPpEt7mTxF77DmbT9pxS4mpngi/LXnQfqYw/Da5WvHOvRqy3b8Bnza
zohuhKK0c4JceJsGbBmrmAJSNSA+bmdPWNnlbxsric3dxIM6B20ojatBeIYa04ah
pM3F4X9+jA2sKStRd9A4vg04cT7tjkK0rBq1rs6aeIBL+Ys62KBrC9HcO98m4IYP
0ZUx04Whl6JQcahhyxj2sEoOw4QaPGVOQ+LH4jbcVqO8BGhCsaxcXrQJEFGy7M4U
yGV/jN58FoAsLR6kCoUgBGhJusl191FqvxYYh5vsUjavznA9iAs5BNvoDH3HgCDy
8Rc7aBvLo02fo0EOPjqXX7SaToRg8/PN3EvfdeiKLlKk3lcIs0FdUAgHmPcWPM3M
+4+mg3js8dFQWYggy5fpsnIk48IWG4AVAq99ElFLEmwxa06CeUsc4MlbpyoM3ySS
ddfIfh6U+WlPFRkOU6Nvz56Kvne3nkGnF0BfkeB3yXHqLvb1IEmEEGUhTRPtv+ai
PX3+8Tmq7mtXXIEew5ypFMHAynnu7qCc7uNMpuzIhLvtuvTc6s7qbci/pm5jCOD6
9eFTz3aVC6gBANyfbjsrvoFt8H1Vh8k/dZXxHXiOdMzDrb+P+grtW8S7X05HFwA3
wUCdQrvSAehLiFqiyFtXibpIxl7+Bop2ClEg43y0AWAt+y6P8cgpBHqmalKhtWxv
6U84KPtSFQqWIzz9r2s9n+GgEQiNSrhPqcelW1j/JFKTy+vnoqbQKu8nTpoxW6Hx
msVL0AQr5+AJU0FeT+LiHx02UlFQPE3iA15klUwpAL11W4bk6oGcPg8jVUlF+5C0
Ny+FCOo0vh3YBSK8FntxHb/7LnAA2UVcqLAXfxQn9rcOqUBG9s0o2iEbRFd1wTMY
0z6pAjy8TkmbLaAHM4ba5x2nAplV2B59wh4XCwbykTsWkCSmiaQW51xbCqqwO63z
kjeAc5P/AdEC5rs4fT1FWOGcAZS0H6fx1rC5QIT6DwEUc0vkQz2wHjFlfXjwGfX8
DmX4mHv0r+xowOQyr25YVewf/W0tC8qAvy9ZsN4P1m9NQ7yuc6jEdzC6T1DUGMpc
JZSZcXwGrEgQn6gBiEof+NKi6+iCCZlcn6mGF/iY3Rcls/uZmtV5k/mQBVwCDfel
u/nY8HAPVZeOzj/xiyUUcESlRHpW6VDSSTr+z/MFAwD+3+MTZVKUGBakGY5nUZY+
r1bO54YQDeyUDdYcigpo2ThjR0VXjO35rBvq2bzBKlPfOHZoxhjqtypKbkyPEp+3
tAJS2ZDy2LYTEYIF5eL/a5kOfIbj9Wjhcav4RMHo3RBXDFgXUF4SZXLp/vTnj658
58jpvfPUBs47rGShFblOqdyfw4rjwAS4y9zA+SFN8vFcnFM+G5SZFXzo9eilTnCR
EOlZr4PaaxJzCh30MfjJMliL3KNlF1A36jBdlghuvoATOdtn5Np83dCvkE8ozPsc
x8Hx7sBloErB11qcMhL1VX0JzbfgIU7bkeQZO+ISF8/ifwfyYjzFHeQbz+F0qziu
5qbXcLD8WEx0xfu9twJcB96xRKBcLvGGT4zbEyCdqCrk567gY5Am1+ozYm1zgvFa
WRg0NhVNQxyXpa5+1S1qLiO3x9YR7xfUVgTKL1PSUU7TyzXJSZNUWTKE8ez7h+e5
OT26gGQrrVgSll1r30oVw2l3KIqJgaYFK0gNQD/iYpRi4UWw5UVFxcjdg8G8xGCd
RxU/y31zWrWYMkWUktwgKHm6dpnoc7OerJwApq7P3TuI/a45DcYONHTH9gV+39S0
ZwFBKJ16E1PzpheD0FQZr6aLzLjwfrlc2ou8EjquwwClCnJVWfHw25XPRni69W2u
LF04ouXT+9jwHbcHIxu7feyTKT45A0wtnubnsxhUqGihOgBg23RLJVWZWmLvwmWs
dQzP40OWG3NqTaNAdGwBYNgiAZ9XSwy17SBy38I1h2EuS1Kqfde6fRz29LXanglB
Y+O3qgC8pmhvx1Q35oo9ENj58iXdsF3Rw+F9q+Uuuv+8dwn2cH5cnrhsjg6fZL/P
CzAET8/7/ZHMyECqkOmPw5Z2CrFp+T1Euhk+uEa5Y8YGQ3bmaKgdPSwxM1m/mTtD
3U/UW7omQP62WVnw2lgYaw0GO6DXzGIt1n6HQJDfaTo36oDAAHonzRGGTjxAqU8U
sIxOsOLG/GOhVUvOMGAk939NXgOlkf2TQ22lsnx+S18mGIeR3xyN08m0SeLPtbEF
QwVd+2leWWewvWE/+Upb9CeTGgSn0IDAmuW1TPAvUdOVEnLCTjMHLPueDOjep+5j
AsABZJreMqvWac3nEm0ZtYvuKiS3GDtGUMQTXW5VPojc/iVqvmZkfdKNywsjh9fp
urKrG7YSGdm+0690BPO9k6LQwWU50AO26229XaeP768tdRjAZt1WtijWN9u3QxkO
tLqCSUf226UPSyFpVXljY8INCOjhUDMS/4cDQalwM8CgmyjNjghG/nD9SdFnIAwd
j9XSHDPZDQww168aRAKcJRQfzcq6q3AU4yXW9He/XhelzGXhMtz89JSNvSFogNbE
XjRg8LI0p1e8/EH6X/Kwde2A4Ov7MZ85Z9B8zxVRMZO3m/rpJQP99WTRlY9KzJTM
xFCLy9oxPgZZYdrwIL281WuHZsXi0OFbt3gRDfHIhvjxIRChV1b4e9yt5RFkRmyL
OHwBEPPXpD3mIPdURoUnbVpIHkRy5IqmV6zIdrqGmOlKuvoo8KNGNsJxsdnP0vxf
ZqZsKUHplfZ95gMcwOX35Je+vpG/iaLb9j2TRQLjrxJBN+0t8HAvxDGAfUpf2ot4
pp1NjCYzwHOKtKB5GlXFz3uH28INYKX3jivbkpYSUt2d9uixPOw21EZv2u8v+OHy
l/vWqG6beDLTRSKrVn3UzDmY4LBpXIYnXEEZ85b/8PSrhVWt82Qn0I1624g7+7Zl
CobrvhGIdEuxedGjeRHG302Jr+J26HtiuMlYdoMd+029tXQ5kdS60Cw6G46G22WW
E/TOiqGyziZTgd1mBAOUwjvWY161v39pP/Z3dCp/UAjAHaVE5GAxlq3EREq8XXNG
rpArUMBbZqJiGH30NTH5FNmhAflBrgKLlMUZMJJ1fJEyj+kUrD1bJFXn6Dh7ADwx
tWs6k5JU96MNUK805TQp5caYQ1NtOrVRqauTD2kz8mJ3RrA4M3b//MqmIBrVkduq
UzbliKVApzcAB8+ZAx7dkez9LAsl0Z1WuWGi/N3CRm0G1Il/eMFARxAp2c+ygnhA
958lWiC/D1MwmD6n9rFYhyxGbAf1TX6bZjLJwxb54ksWiiaPL5YANNKSMfeiR2am
rrOEJL35oCQZqFige/nuvbnWtSMjEVqFrC4xmESvU4V78RbxkBWAhDJQUG5Oy4XW
N3Vq9P4YwBCHX4eqvDofUo8DUHRyLKZ9fIOMqTT93iUT13QLik/EEWFgcA1V03Xd
BY8hRSXK1GCYkL84sZ+9ThMhPcDcvtMuF6Vf5XxtOR2Xd++574vAPoWOZpZKv4uA
AvgY2wvDrhmjosSfHk7C7eJLvQChcAd+nlAq8F5xoRNdf7f2jWdBQdiNJX3zQ8kg
lZWHeBiwRuzjOw7nEf7Ul+4+D2AE2QK1KLCNkJd7I/Uuq2KH/hrS8clyTZ5MGB5M
TdZxOAULeHDb5j2HS8+owrjsfuoNPzzaeJ8NALcaULcmuUaCOEeYlFlb9dMgf+ar
9kTt2fe3qYzP3rPm1cCbb18u3dEdtSaSTd+pNJTKZ726ud/K2uzBh6IPKMUXF992
07SODSEffcxBmDcKn3L+B8dSyl9P8OyCmk0sCt9Jw6R31xILzJySiE3OZgI+8LdJ
MvI4f1xcPVZO39zacqBrDQOZG+koVvG5shlo8zj/2ou3uGtTLbn5cBCLHYN/ec6h
5Z9aZxcEJhODKF4b0UoK7sDnXtI0oj1gUilFMyF4pNdwypfrzqG1MpWFLGS3OxgV
pN//xgx3K4RynvDbU2tbj36c/X9z1T48OftdtsGCu1hmimRxKJ0jImlEJ7DDWar1
P9iB8FziWC8q/bphIIqpjBO+AtOuF2SQU3RYw54viex41/a6wfI5c8qUyLDsJfuc
vLF5OY2KNudjFiZfxrbFyt1t0xFPWXaWb3JJiPMTY9QCF32u5zN0NsK8+Aw/lNaT
Xwrr3CVcDbLM3On7u0lMUxdy1H8Fd+P7xFxjC0ArhHtgPwDvO42PcfUKpkYGBWwo
cCwn4JprQKbCyCN2/doKLlVvZKTE86WYdmLIGGP08FxAkPhT6gNa6U7GEOasbjmm
dMKc+zkadGbbfYq5ks/k5DGj4oIoXof4MzXhURRz5kUQL/knN/L+2FW3zMWb/8GW
oCOKKcwMvz0fTyUhYJQH1n8ovwq4ilQGNhk4tTAdwk8=
`protect END_PROTECTED
