///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company:			
//				
// Engineer:		
//
// Create Date:		
// Design Name:		
// Module Name:		
// Project Name:	
// Target Devices:  
// Tool versions:
// Description:		
//
// Dependencies:
//	 
// 	 
//
// Revision:
//
//
//
//
// Additional Comments:     
//                          
//                          
//                          
//                          
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`ifndef __CNN_LAYER_ACCEL_AWP__
`define __CNN_LAYER_ACCEL_AWP__


//---------------------------------------------------------------------------------------------------------------------------------------------------
// Includes
//---------------------------------------------------------------------------------------------------------------------------------------------------
`include "utilities.svh"


`define CONVMAP_FIFO_WR_WTH                	1024 // TODO: Remove hard coding
`define CONVMAP_FIFO_RD_WTH                	1024 // TODO: Remove hard coding
`define CONVMAP_FIFO_RD_DTH					512	 // TODO: Remove hard coding
`define MAX_AWPS                            1

`endif