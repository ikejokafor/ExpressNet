`ifndef	__CNL_SC2_GENERATOR__
`define	__CNL_SC2_GENERATOR__


`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company:			
//				
// Engineer:		
//
// Create Date:		
// Design Name:		
// Module Name:		
// Project Name:	
// Target Devices:  
// Tool versions:
// Description:		
//
// Dependencies:
//	 
// 	 
//
// Revision:
//
//
//
//
// Additional Comments:     This class creates test for DUT
//                              pre_randomize() and post_randomize() are built in overridable functions  
//                          Not testing padding > 1
//                          
//                          floor((W - F + (2 * P)) / S) + 1
//                          
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`include "cnn_layer_accel.svh"
`include "cnn_layer_accel_AWP.svh"
`include "cnn_layer_accel_conv1x1_pip.svh"
`include "cnn_layer_accel_FAS.svh"
`include "cnn_layer_accel_FAS_pip_ctrl.svh"
`include "cnn_layer_accel_QUAD.svh"
`include "cnn_layer_accel_trans_fifo.svh"
`include "awe.svh"
`include "axi_defs.svh"

`include "generator.sv"
`include "cnl_sc2_verif_defs.svh"
`include "cnn_layer_accel_verif_defs.svh"


class `scX_genParams_t extends genParams_t;
endclass: `scX_genParams_t


class `scX_crtTestParams_t extends crtTestParams_t;
    int num_input_rows;
    int num_input_cols;
    int depth;
    int num_kernels;
    int stride;
    int padding;
    int kernel_size;
    int conv_out_fmt;
    bool upsample;
    int cascade;
endclass: `scX_crtTestParams_t


class `cnl_scX_generator extends generator;
    extern function new(genParams_t genParams = null);
    extern function void createTest(crtTestParams_t params);
    extern function void plain2bits();
    extern function void post_randomize();
    

    rand int m_num_input_rows                                                           ;
    rand int m_num_input_cols                                                           ;
    int      m_num_expd_input_cols                                                      ;
    int      m_num_expd_input_rows                                                      ;
    int      m_num_input_rows_cfg                                                       ;
    int      m_num_input_cols_cfg                                                       ;
    int      m_num_output_rows_cfg                                                      ;
    int      m_num_output_cols_cfg                                                      ;
    int      m_num_output_rows                                                          ;
    int      m_num_output_cols                                                          ;    
    int      m_num_acl_output_rows                                                      ;
    int      m_num_acl_output_cols                                                      ;
    int      m_pfb_full_count_cfg                                                       ;
    rand int m_depth                                                                    ;
    rand int m_num_kernels                                                              ;
    rand int m_kernel_size                                                              ;
    rand int m_stride                                                                   ;
    rand int m_padding                                                                  ;
    int m_uple_fctr                                                                     ;
    bool m_upsample                                                                     ;
    int m_conv_out_fmt                                                                  ;
    int m_num_expd_input_cols_cfg                                                       ;
    int m_num_expd_input_rows_cfg                                                       ;
    int m_crpd_input_col_start_cfg                                                      ;
    int m_crpd_input_row_start_cfg                                                      ;
    int m_crpd_input_col_end_cfg                                                        ;
    int m_crpd_input_row_end_cfg                                                        ;
    int m_pix_seq_data_full_count_cfg                                                   ;
    int m_cascade_cfg                                                                   ;
    int m_num_kernels_cfg                                                               ;
    int m_pix_data[]                                                                    ;
    int m_pix_data_upsle[]                                                              ;
    int m_kernel_data[]                                                                 ;
    logic [15:0] m_pix_seq_data_sim[0:((`MAX_NUM_INPUT_COLS * `NUM_CE_PER_QUAD) - 1)]   ;
    logic [15:0] m_pix_data_sim[]                                                       ;
    logic [15:0] m_pix_data_upsle_sim[]                                                 ;
    logic [15:0] m_kernel_data_sim[]                                                    ;
    

    constraint c0 {      
        solve m_num_input_rows before m_num_input_cols;
        m_num_input_rows inside {[`MIN_NUM_INPUT_ROWS:`MAX_NUM_INPUT_ROWS]};
        m_num_input_cols == m_num_input_rows;
        m_depth == `NUM_CE_PER_QUAD;
        m_kernel_size == 3;
        m_num_kernels inside {[1:`MAX_BRAM_3x3_KERNELS]};
        m_stride inside {[1:2]};
        m_padding inside {[0:`MAX_PADDING]};
        m_upsample inside {[0:1]};
    }
endclass: `cnl_scX_generator


function `cnl_scX_generator::new(genParams_t genParams = null);
    `scX_genParams_t `scX_genParams;


    if(genParams != null) begin
        $cast(`scX_genParams, genParams);
        m_ti = `scX_genParams.ti;
        m_outputDir = `scX_genParams.outputDir;
    end
endfunction: new


function void `cnl_scX_generator::createTest(crtTestParams_t params);
    `scX_crtTestParams_t `scX_crtTestParams;
    
    
    $cast(`scX_crtTestParams, params);
    m_num_input_rows = `scX_crtTestParams.num_input_rows;
    m_num_input_cols = `scX_crtTestParams.num_input_cols;
    m_depth = `scX_crtTestParams.depth;
    m_num_kernels = `scX_crtTestParams.num_kernels;
    m_kernel_size = `scX_crtTestParams.kernel_size;
    m_conv_out_fmt = `scX_crtTestParams.conv_out_fmt;
    m_stride = `scX_crtTestParams.stride;
    m_padding = `scX_crtTestParams.padding;
    m_upsample = `scX_crtTestParams.upsample;
    m_cascade_cfg = `scX_crtTestParams.cascade;
    post_randomize();

    
    $display("// Created Specific Test ----------------------------------------");
    $display("// Test Index:            %0d", m_ti                              );
    $display("// Num Input Rows:        %0d", m_num_input_rows                  );
    $display("// Num Input Cols:        %0d", m_num_input_cols                  );
    $display("// Input Depth:           %0d", m_depth                           );
    $display("// Num Kernels:           %0d", m_num_kernels                     );
    $display("// Kernel size:           %0d", m_kernel_size                     );
    $display("// Stride                 %0d", m_stride                          );
    $display("// Padding:               %0d", m_padding                         );
    $display("// Upsample               %0d", m_upsample                        );
    $display("// Num Output Rows:       %0d", m_num_output_rows                 );
    $display("// Num Output Cols:       %0d", m_num_output_cols                 );
    $display("// Num Acl Output Rows:   %0d", m_num_acl_output_rows             );
    $display("// Num Acl Output Cols:   %0d", m_num_acl_output_cols             );
    $display("// Conv Output Format:    %0d", m_conv_out_fmt                    );
    $display("// Created Specific Test ----------------------------------------");
    $display("\n");

endfunction: createTest


function void `cnl_scX_generator::plain2bits();
    int i;
    int j;
    int a;
    int b;
    int n;


    m_pix_data_sim = new[m_pix_data.size()];
    foreach(m_pix_data[i]) begin
        m_pix_data_sim[i] = m_pix_data[i];
    end

    
    if(m_upsample) begin
        m_pix_data_upsle_sim = new[m_pix_data_upsle.size()];
        foreach(m_pix_data_upsle[i]) begin
            m_pix_data_upsle_sim[i] = m_pix_data_upsle[i];
        end
    end
    
    
    m_kernel_data_sim = new[m_num_kernels * m_depth * `KERNEL_3x3_COUNT_FULL];
    for(i = 0; i < m_num_kernels; i = i + 1) begin
        for(j = 0; j < m_depth; j = j + 1) begin
            n = 0;
            for(a = 0; a < m_kernel_size; a = a + 1) begin
                for(b = 0; b < m_kernel_size; b = b + 1) begin
                    m_kernel_data_sim[(i * m_depth + j) * `KERNEL_3x3_COUNT_FULL + n]
                        = m_kernel_data[((i * m_depth + j) * m_kernel_size + a) * m_kernel_size + b];
                    n = n + 1;
                end
            end
            m_kernel_data_sim[(i * m_depth + j) * `KERNEL_3x3_COUNT_FULL + n] = 0;
        end
    end
endfunction: plain2bits


function void `cnl_scX_generator::post_randomize();
    int i;
    int j;
    int k;
    int a;
    int b;
    shortreal fl_num_expd_input_rows;
    shortreal fl_num_expd_input_cols;
    shortreal fl_num_input_cols;
    int fl_pix_seq_data_full_count;
    int in_index;
    int out_index;
    int num_conv_input_rows;
    int num_conv_input_cols;


    m_depth = m_depth * `NUM_QUADS;
    m_num_kernels_cfg = m_num_kernels - 1;
    m_num_output_rows = ((m_num_input_rows - m_kernel_size + (2 * m_padding)) / m_stride) + 1;
    m_num_output_cols = ((m_num_input_rows - m_kernel_size + (2 * m_padding)) / m_stride) + 1;     
    if(m_padding && !m_upsample) begin
        m_num_expd_input_rows = m_num_input_rows + 2;
        m_num_expd_input_cols = m_num_input_cols + 2;       
    end else if(!m_padding && m_upsample) begin
        m_num_expd_input_rows = m_num_input_rows * 2;
        m_num_expd_input_cols = m_num_input_cols * 2; 
        m_num_output_rows = ((m_num_expd_input_rows - m_kernel_size + (2 * m_padding)) / m_stride) + 1;
        m_num_output_cols = ((m_num_expd_input_cols - m_kernel_size + (2 * m_padding)) / m_stride) + 1;
    end else if(m_padding && m_upsample) begin
        m_num_expd_input_rows = (m_num_input_rows * 2) + 2;
        m_num_expd_input_cols = (m_num_input_cols * 2) + 2;
        m_num_output_rows = (((m_num_expd_input_rows - 2) - m_kernel_size + (2 * m_padding)) / m_stride) + 1;
        m_num_output_cols = (((m_num_expd_input_cols - 2) - m_kernel_size + (2 * m_padding)) / m_stride) + 1;        
    end else begin // !m_padding && !m_upsample
        m_num_expd_input_rows = m_num_input_rows;
        m_num_expd_input_cols = m_num_input_cols;      
    end
    m_num_input_rows_cfg                = m_num_input_rows - 1;
    m_num_input_cols_cfg                = m_num_input_cols - 1;   
    m_num_expd_input_rows_cfg           = m_num_expd_input_rows - 1;
    m_num_expd_input_cols_cfg           = m_num_expd_input_cols - 1;      
    m_crpd_input_col_start_cfg          = 1;
    m_crpd_input_row_start_cfg          = 1;
    m_crpd_input_row_end_cfg            = m_num_expd_input_rows - 2;
    m_crpd_input_col_end_cfg            = m_num_expd_input_cols - 2;
    m_pfb_full_count_cfg                = m_num_expd_input_cols;
    

    if(m_padding && m_stride == 2) begin    
        fl_num_expd_input_rows          = m_num_expd_input_rows;
        fl_num_expd_input_cols          = m_num_expd_input_cols;
        m_num_acl_output_rows           = $ceil(fl_num_expd_input_rows / shortreal'(2)) - 1;
        m_num_acl_output_cols           = $ceil(fl_num_expd_input_cols / shortreal'(2));
        m_num_output_rows_cfg           = $ceil(fl_num_expd_input_rows / shortreal'(2)) - 1;
        m_num_output_cols_cfg           = $ceil(fl_num_expd_input_cols / shortreal'(2));
        m_pix_seq_data_full_count_cfg   = `WINDOW_3x3_NUM_CYCLES * $ceil(fl_num_expd_input_cols / shortreal'(2));
    end else if(!m_padding && m_stride == 2) begin
        fl_num_expd_input_rows          = m_num_expd_input_rows;
        fl_num_expd_input_cols          = m_num_expd_input_cols;
        m_num_acl_output_rows           = $ceil(fl_num_expd_input_rows / shortreal'(2)) - 1;
        m_num_acl_output_cols           = $ceil(fl_num_expd_input_cols / shortreal'(2));
        m_num_output_rows_cfg           = $ceil(fl_num_expd_input_rows / shortreal'(2)) - 1;
        m_num_output_cols_cfg           = $ceil(fl_num_expd_input_cols / shortreal'(2));
        m_pix_seq_data_full_count_cfg   = `WINDOW_3x3_NUM_CYCLES * $ceil(fl_num_expd_input_cols / shortreal'(2)); 
    end else if(m_padding && m_stride == 1) begin
        m_num_acl_output_rows           = (((m_num_expd_input_rows - 2) - m_kernel_size + (2 * m_padding)) / m_stride) + 1;
        m_num_acl_output_cols           = m_num_expd_input_cols;
        m_num_output_rows_cfg           = (((m_num_expd_input_rows - 2) - m_kernel_size + (2 * m_padding)) / m_stride) + 1;
        m_num_output_cols_cfg           = m_num_expd_input_cols;
        m_pix_seq_data_full_count_cfg   = `WINDOW_3x3_NUM_CYCLES * m_num_expd_input_cols;
    end else begin // (!m_padding && m_stride == 1)
        m_num_acl_output_rows           = ((m_num_expd_input_rows - m_kernel_size + (2 * m_padding)) / m_stride) + 1;
        m_num_acl_output_cols           = m_num_expd_input_cols;
        m_num_output_rows_cfg           = ((m_num_expd_input_rows - m_kernel_size + (2 * m_padding)) / m_stride) + 1;
        m_num_output_cols_cfg           = m_num_expd_input_cols;
        m_pix_seq_data_full_count_cfg   = `WINDOW_3x3_NUM_CYCLES * m_num_expd_input_cols;
    end


    m_pix_data = new[m_depth * m_num_input_rows * m_num_input_cols];
    foreach(m_pix_data[i]) begin
        m_pix_data[i] = $urandom_range(`MIN_RND_VALUE, `MAX_RND_VALUE);
    end
    

    if(m_upsample) begin
        m_uple_fctr = 2;
        if(m_padding) begin
            num_conv_input_rows = m_num_expd_input_rows - 2;
            num_conv_input_cols = m_num_expd_input_cols - 2;
        end else begin
            num_conv_input_rows = m_num_expd_input_rows;
            num_conv_input_cols = m_num_expd_input_cols;
        end
        m_pix_data_upsle = new[m_depth * num_conv_input_rows * num_conv_input_cols]; 
        for(k = 0; k < m_depth; k = k + 1) begin
            for(j = 0; j < m_num_input_rows * m_uple_fctr; j = j + 1) begin
                for(i = 0; i < m_num_input_cols * m_uple_fctr; i = i + 1) begin
                    in_index = k * m_num_input_cols * m_num_input_rows + (j / m_uple_fctr) * m_num_input_cols + i / m_uple_fctr;
                    out_index = k * m_num_input_cols * m_num_input_rows * m_uple_fctr * m_uple_fctr + j * m_num_input_cols * m_uple_fctr + i;
                    m_pix_data_upsle[out_index] = m_pix_data[in_index];
                end
            end
        end
    end
 

    m_kernel_data = new[m_num_kernels * m_depth * m_kernel_size * m_kernel_size]; 
    for(i = 0; i < m_num_kernels; i = i + 1) begin
        for(j = 0; j < m_depth; j = j + 1) begin
            for(a = 0; a < m_kernel_size; a = a + 1) begin
                for(b = 0; b < m_kernel_size; b = b + 1) begin
                    m_kernel_data[((i * m_depth + j) * m_kernel_size + a) * m_kernel_size + b] = $urandom_range(`MIN_RND_VALUE, `MAX_RND_VALUE);
                end
            end
        end
    end
    
 
    // BEGIN logic ----------------------------------------------------------------------------------------------------------------------------------
    if(m_stride == 1) begin
        // RM = Row matriculate
        // RST = Reset MACC reg
        // P = parity bit
        // SEQ = sequence value
        //
        //                             RM    RST   P     SEQ
        m_pix_seq_data_sim[0] = {3'b0, 1'b0, 1'b1, 1'b1, 10'd0  };
        m_pix_seq_data_sim[1] = {3'b0, 1'b0, 1'b0, 1'b0, 10'd2  };
        m_pix_seq_data_sim[2] = {3'b1, 1'b0, 1'b0, 1'b0, 10'd512};
        m_pix_seq_data_sim[3] = {3'b0, 1'b0, 1'b0, 1'b0, 10'd513};
        m_pix_seq_data_sim[4] = {3'b0, 1'b1, 1'b0, 1'b0, 10'd514};

        j = 0;
        for(i = `WINDOW_3x3_NUM_CYCLES; i < (`MAX_NUM_INPUT_COLS * `WINDOW_3x3_NUM_CYCLES); i = i + `WINDOW_3x3_NUM_CYCLES) begin            
            if((j % 2) == 0) begin
                m_pix_seq_data_sim[i    ] = {3'b0, 1'b0, 1'b1, 1'b0, m_pix_seq_data_sim[i - 5][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd1};
                m_pix_seq_data_sim[i + 1] = {3'b0, 1'b0, 1'b0, 1'b1, m_pix_seq_data_sim[i - 4][`PIX_SEQ_DATA_SEQ_FIELD]};
            end else begin           
                m_pix_seq_data_sim[i    ] = {3'b0, 1'b0, 1'b1, 1'b1, m_pix_seq_data_sim[i - 5][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd1};
                m_pix_seq_data_sim[i + 1] = {3'b0, 1'b0, 1'b0, 1'b0, m_pix_seq_data_sim[i - 4][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd2};
            end
            m_pix_seq_data_sim[i + 2] = {3'b1, 1'b0, 1'b0, 1'b0, m_pix_seq_data_sim[i - 3][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd1};
            m_pix_seq_data_sim[i + 3] = {3'b0, 1'b0, 1'b0, 1'b0, m_pix_seq_data_sim[i - 2][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd1};
            m_pix_seq_data_sim[i + 4] = {3'b0, 1'b1, 1'b0, 1'b0, m_pix_seq_data_sim[i - 1][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd1};
            j = (j + 1) % 2;
        end
        while(i < (`MAX_NUM_INPUT_COLS * `NUM_CE_PER_QUAD)) begin
            m_pix_seq_data_sim[i] = 0;
            i = i + 1;
        end
    end else if(m_stride == 2) begin
        // RM = Row matriculate
        // RST = Reset MACC reg
        // P = parity bit
        //                            RM   RST    P
        m_pix_seq_data_sim[0] = {3'b0, 1'b0, 1'b1, 1'b1, 10'd0  };
        m_pix_seq_data_sim[1] = {3'b0, 1'b0, 1'b0, 1'b0, 10'd2  };
        m_pix_seq_data_sim[2] = {3'b1, 1'b0, 1'b0, 1'b0, 10'd512};
        m_pix_seq_data_sim[3] = {3'b1, 1'b1, 1'b0, 1'b0, 10'd513};
        m_pix_seq_data_sim[4] = {3'b0, 1'b1, 1'b0, 1'b0, 10'd514};
    
        j = 0;
        for(i = `WINDOW_3x3_NUM_CYCLES; i < ((`MAX_NUM_INPUT_COLS / 2) * `WINDOW_3x3_NUM_CYCLES); i = i + `WINDOW_3x3_NUM_CYCLES) begin
            m_pix_seq_data_sim[i    ] = {3'b0, 1'b0, 1'b1, 1'b1, m_pix_seq_data_sim[i - 5][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd2};
            m_pix_seq_data_sim[i + 1] = {3'b0, 1'b0, 1'b0, 1'b0, m_pix_seq_data_sim[i - 4][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd2};
            m_pix_seq_data_sim[i + 2] = {3'b1, 1'b0, 1'b0, 1'b0, m_pix_seq_data_sim[i - 3][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd2};
            m_pix_seq_data_sim[i + 3] = {3'b1, 1'b1, 1'b0, 1'b0, m_pix_seq_data_sim[i - 2][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd2};
            m_pix_seq_data_sim[i + 4] = {3'b0, 1'b1, 1'b0, 1'b0, m_pix_seq_data_sim[i - 1][`PIX_SEQ_DATA_SEQ_FIELD] + 10'd2};
            j = (j + 1) % 2;
        end
        while(i < (`MAX_NUM_INPUT_COLS * `NUM_CE_PER_QUAD)) begin
            m_pix_seq_data_sim[i] = 0;
            i = i + 1;
        end
    end
    // END logic ------------------------------------------------------------------------------------------------------------------------------------

endfunction: post_randomize


`endif