`ifndef __CNL_SC1_VERIF_DEFS__
`define __CNL_SC1_VERIF_DEFS__


`define cnl_scX_DUTOutput       cnl_sc1_DUTOutput
`define cnl_scX_generator       cnl_sc1_generator
`define cnl_scX_monitor         cnl_sc1_monitor
`define cnl_scX_scoreboard      cnl_sc1_scoreboard
`define cnl_scX_agent           cnl_sc1_agent
`define cnl_scX_assertion       cnl_sc1_assertion
`define cnl_scX_driver          cnl_sc1_driver
`define cnl_scX_environment     cnl_sc1_environment

`define scX_DUTOutParams_t      sc1_DUTOutParams_t
`define scX_datum_t             sc1_datum_t
`define scX_genParams_t         sc1_genParams_tarams_t
`define scX_crtTestParams_t     sc1_crtTestParams_t
`define scX_monParams_t         sc1_monParams_t
`define scX_scoreParams_t       sc1_scoreParams_t
`define scX_agentParams_t       sc1_agentParams_t
`define scX_asrtParams_t        sc1_asrtParams_t
`define scX_drvParams_t         sc1_drvParams_t


`define scX_DUTOutParams        sc1_DUTOutParams
`define scX_datum               sc1_datum
`define scX_genParams           sc1_genParams_tarams
`define scX_crtTestParams       sc1_crtTestParams
`define scX_monParams           sc1_monParams
`define scX_scoreParams         sc1_scoreParams
`define scX_agentParams         sc1_agentParams
`define scX_asrtParams          sc1_asrtParams
`define scX_drvParams           sc1_drvParams
`define scX_query               sc1_query
`define scX_test                sc1_test
`define scX_sol                 sc1_sol


`endif
