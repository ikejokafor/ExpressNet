library verilog;
use verilog.vl_types.all;
entity cnn_layer_accel_quad_intf is
    port(
        clk_if          : in     vl_logic;
        clk_core        : in     vl_logic;
        rst             : out    vl_logic;
        job_start       : out    vl_logic;
        job_accept      : in     vl_logic;
        job_parameters  : out    vl_logic_vector(127 downto 0);
        job_fetch_request: in     vl_logic;
        job_fetch_ack   : out    vl_logic;
        job_fetch_complete: out    vl_logic;
        job_complete    : in     vl_logic;
        job_complete_ack: out    vl_logic;
        cascade_in_valid: out    vl_logic;
        cascade_in_ready: in     vl_logic;
        cascade_in_data : out    vl_logic_vector(127 downto 0);
        cascade_out_valid: in     vl_logic;
        cascade_out_ready: out    vl_logic;
        cascade_out_data: in     vl_logic_vector(127 downto 0);
        config_valid    : out    vl_logic_vector(3 downto 0);
        config_accept   : in     vl_logic_vector(3 downto 0);
        config_data     : out    vl_logic_vector(127 downto 0);
        weight_valid    : out    vl_logic;
        weight_ready    : in     vl_logic;
        weight_data     : out    vl_logic_vector(127 downto 0);
        result_valid    : in     vl_logic;
        result_accept   : out    vl_logic;
        result_data     : in     vl_logic_vector(15 downto 0);
        pixel_valid     : out    vl_logic;
        pixel_ready     : in     vl_logic;
        pixel_data      : out    vl_logic_vector(127 downto 0);
        num_input_cols_cfg: out    vl_logic_vector(9 downto 0);
        num_input_rows_cfg: out    vl_logic_vector(9 downto 0);
        pfb_full_count_cfg: out    vl_logic_vector(9 downto 0);
        kernel_full_count_cfg: out    vl_logic_vector(7 downto 0);
        kernel_group_cfg: out    vl_logic_vector(6 downto 0);
        convolution_stride_cfg: out    vl_logic_vector(6 downto 0);
        kernel_size_cfg : out    vl_logic_vector(4 downto 0);
        padding_cfg     : out    vl_logic_vector(4 downto 0);
        upsample_cfg    : out    vl_logic;
        num_kernel_cfg  : out    vl_logic_vector(6 downto 0);
        num_output_rows_cfg: out    vl_logic_vector(9 downto 0);
        num_output_cols_cfg: out    vl_logic_vector(9 downto 0);
        pix_seq_data_full_count_cfg: out    vl_logic_vector(11 downto 0);
        pded_num_input_cols_cfg: out    vl_logic_vector;
        pded_num_input_rows_cfg: out    vl_logic_vector;
        crpd_input_col_start_cfg: out    vl_logic_vector;
        crpd_input_row_start_cfg: out    vl_logic_vector;
        crpd_input_col_end_cfg: out    vl_logic_vector;
        crpd_input_row_end_cfg: out    vl_logic_vector;
        output_row      : in     integer;
        output_col      : in     integer;
        output_depth    : in     integer
    );
end cnn_layer_accel_quad_intf;
