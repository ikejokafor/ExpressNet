`ifndef __CNL_SC0_VERIF_DEFS__
`define __CNL_SC0_VERIF_DEFS__


`define cnl_scX_DUTOutput       cnl_sc0_DUTOutput
`define cnl_scX_generator       cnl_sc0_generator
`define cnl_scX_monitor         cnl_sc0_monitor
`define cnl_scX_scoreboard      cnl_sc0_scoreboard
`define cnl_scX_agent           cnl_sc0_agent
`define cnl_scX_assertion       cnl_sc0_assertion
`define cnl_scX_driver          cnl_sc0_driver
`define cnl_scX_environment     cnl_sc0_environment

`define scX_DUTOutParams_t      sc0_DUTOutParams_t
`define scX_datum_t             sc0_datum_t
`define scX_genParams_t         sc0_genParams_tarams_t
`define scX_crtTestParams_t     sc0_crtTestParams_t
`define scX_monParams_t         sc0_monParams_t
`define scX_scoreParams_t       sc0_scoreParams_t
`define scX_agentParams_t       sc0_agentParams_t
`define scX_asrtParams_t        sc0_asrtParams_t
`define scX_drvParams_t         sc0_drvParams_t


`define scX_DUTOutParams        sc0_DUTOutParams
`define scX_datum               sc0_datum
`define scX_genParams           sc0_genParams_tarams
`define scX_crtTestParams       sc0_crtTestParams
`define scX_monParams           sc0_monParams
`define scX_scoreParams         sc0_scoreParams
`define scX_agentParams         sc0_agentParams
`define scX_asrtParams          sc0_asrtParams
`define scX_drvParams           sc0_drvParams
`define scX_query               sc0_query
`define scX_test                sc0_test
`define scX_sol                 sc0_sol


`endif
