`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgqZw9iLAr8AyzA3J9O9SgSo5VA4Lvi0EbJn11fdYGLVb8C28Q4581jTG/jPQNIU
RBJwDYOQfPZvKvrgfHyrWabpWniJUrKV3vSIEsjgsNFmW5YNSIAH6YCnc7xunafy
Gy4/QS/ismHpTHHUdGmJBziluJttettcS7N7qL3qe6aIypwbHaC+7xifPPktXvXY
q/EqZFtYl89SxqbulGd4Zr5ZcoeNvO1PRmjBfM9gDIisWMbuYHtASb2XCzUi0v8S
Kt4ZEq2gtZ7dTRyTWj1y1LxgYSYGx4305ZcW6osn+Aqq1BjN1mg9cLUvynXvsUX3
bSZmGJss4AzEJODfkq8xHYK9D9Ihu5Q5N1wL41fujjClzIvWG4ntDt0MFKiSlDx9
OOXEhMaEvkGRpNiO4dTVP7qmnearsWlnkSIA4lzLQe7PBLcj3ywa1lcQbwJD0CAJ
aIkx4SSn1OeIlOgMfvQdIPaqs/L1oQpgOGIVUCq9OF2Bf30iVYyayWCibDUc2c1W
QgW/tatSKl6LKV1mvGDkJqae7QMWiW5c3PQnj9EMFuVubGaLdbsvI9dKCX6UujGi
5WzSg0h905gU23qHtaFRydrjeda0OqdIN0bwaKgnLoDquwJAzyW9VYJk2MrW4uFi
/5Qu4TVlvaJFFv46RpWgH6voCgIZwW0cUFQMHJrYRuxP3Fi/weAQSb1y5RXXGagH
6PlcIEJ7qblP75Xx4I1VKq9Bxe/MLtnsaEmhCl1RBdFRGQCLImEmrd68unySDGrU
OS56koCc2M+bGxUm2oMN19Ty6fDH4Vu1xdFKud4yaN5BwD9Brjd69pOA8sdTs+2w
5q1umwNMQswIUTflxpC6kPWziaRpf3LxFWoFNI1pXUzsSO4Eze8H4cNACjniILfB
9AJkEEHGUv0q1TUdBpFjW6oSjlbp7JfKFA6pdSbWcXp8FmqzXJgy1hFHuUriEV/h
e9+0cgqMK4fPZsKJS1BVcikwG1hieih65NM+mrwxaIYz9IxwGFQHVPo93ZkSHwa5
oMg8tITFFMxjxXUdFSW/HqprqxE45wMdwiyFXrmkCY4GtONo7dN8gIeBDDqIug6t
AKfRHpWp091k7LYvm1ZFTpgXnZkcwLdhKcTgu5nJFKtxAxSJM+v8XMId1rFofmu8
iiL1dqk2tOH/SLdH5swQeJrdwN7XustGcj8whTv/Jq9LJjYIsxBwzgAeUshxy8G3
xbAcNt1l7LqQedmPTtUhel9uy37cVNVsGFY0bd+SE/Kj6MNnxOXsPjp9iaxaYEav
BHyLuXbM1GxHMdmYueAcpLyiD1nWQ9JepjjE77PPRwV2GyiggjG9ZIl4tVAMjXZD
6AebNoV9wBT+H2sbIu4Pq97Z7zWqoFvgFErDiq5KDN1XCJa5fFYNluwXrnXDkMMz
w7Xi0uFi1cUddtUEnMkpkHYDGRRVWXeG53ltEWW+pzLPeWQdU85qiZuktPCcqsk4
3UOJMrOqXGbOOqu9/zyQmz26O/zL+uEb++HLjzAnTso7QsKeW0IIsigqsMPWyiyQ
qe0cfCf1TuOZkWRxige58NG4cj+XvctfrAOwbyMeNVaxwcKlMCQ19uGxhpxP8Q39
+GsXi3HIguzW4CwPp7v2StHJcDvSVWxsip+LInmzCPJgQ3g6QzPUuANCKTFv++wB
5/f8EPIbKM9kDm6bDY5VOZRMs4eNthXZ29CY6Kg+wOujcOZZEk6sYsBwXvV3o3sV
UAAaEbuDJeeh5F2Q2S2l6wd0nDVyDAAZ8M5vMIY5Im8KwYUMg7Z8gu1aLR3V3Fj8
8Ll7noho5tuE31mXzYRGYKOhMXc1SXufTloNIL35RwwZL/j2CdMY4mtCGn9Yb++Z
qtS0trAtmZ2P5EXy04kOYEFIlAg16Gipbtx5NL34Kn0D1nB3bDiGMth3RVCcjWgy
iIBnAYzk76qB6nfHuZ+Ojr1fuG65vFpxEMWjRNN9Eveqdv2i7Y7tu8WBeb71sZFD
Ge2mrVk7dqT4o7gHauBl3VfYEm/YKQC6TXRFSPDj2ZlPKH3X9Xv95cbPxzZgGsjM
MPhzTZq/e6YM4YnDFD0YcQIMEYeD6W8KiYgmakOwgWAY1RYJWt79LPgJj2bLEdco
fGLJdgwJoNetPAouDNVmpUKMqhZmkz4OUzEMGIYlW8EuDdjtXR37gWn6io69Sfri
LYK8lcejh/c/6w638wjkq6lazXx5mSEegBjEGAcWOr1NM/8Xz3JOwadRWlexbaVt
RGhxYtogwSvIE2L1TZyoW/0DOdsj4oofyNDP98yCEsjS9+AzKbIdn7v1pT+pKRKi
ngWQTXooCaIv5JPHn8bgOjFykYVRdUvlzee1ozi/uwPXY4kNilu27VtkbT+L6BhX
2BYaTxcQlItF+WFm/7x8y7vdM+CzQMr+AHZsyol4o8Vn+3M+WnbK2+tm/KtK+oX1
q3aLPyrgxE8e0CoQ6HxvbqZcLyU8pQVkHznZfymN+pNfMvArHNTzTsZjq1lQZsuv
GNAbmETKX2QFYR/SPe733vOa13RbwbCD0Ow6rcEbo0RC5E8+ogR/3byXu/PnxAY3
oZgksjcSFEF/ZxLT6MnepF1uIMCilifQpyQUJJP7ujgZNTB7WcWkOBQmwYnyvBBA
kixhEeI8mYbvvdGAROXhjlHbW/II/P97rlCFYVPWVuqQzi2RagfmTZY09v0rv/bt
my7/Bc+4Sh2JvU+hPKtBXwhznNcHfpgno123lCPxGqQYA2iaqCH2fQnLiE6YmA+R
d1CqOAbk3npmyOrtX3aVAJgUPfHM5Ovl4JCQ0rE0p55BILKh2DswM1n+JMf+UFb4
lun66NgK7D9aJGhpdsaplVrf3Tup6aDbKPsJV/BQ3+hNGZAJcmli2v2tuCOi8mSe
zSkS1slPRtvnqdbL15l12h2Lz6SpA3cCH0bJ5S6dRntlYZg5oMdlbvsAB1DcURyL
5qWE69seumHVGFV140oSVbL7faZuIGFU+BMax96zevTDRxV2ZhARyCzQB8qsQbjp
bqeSQt6nhvJ1a8DtGgpWWTqr4Y4FsHZQLZtrIRUfWk08O1YugCElJVjH1tCrJ25a
wMbogqIFzsgwIvDy6+YrZN5yw+KomKAXgPdmFMRvF6ygF1jUINUzVecVzSt10DX4
uUVR3KyCh5VCrAsNzMSBqYD5R4rtBlDKRmwrtSUlwJU3cSPAXlvAD2UxbSQcaiVK
NQ3UPJ5TzE/HUNeHA2xoSiErVGkV00nrjB0Rq3H/hImKKRaQOC8wdBXetrpWmskA
oSbjLXc/1T0zr52s+uTWCfsQ/rGLsE+uvc7e4qjKw1OvDAZYupuqOxb3aux/Jaf+
1/yMcXBPdbM2S85r4UAcf/jt4cMfCENAw/lY/t4856GJ6ufbNwtJmURGwpQ0H7js
mDQd7ZodwYAG854lE/cVXPraHaf6ENG58dIvS3hhlXTgsYgizyGNJhDeqVl4ovXM
YB68H8/9nbAW25AwkVQs4CNY8+dr6SRHJD5MWsEozAgFJ3sUMvShT5I/uUDzNENH
PQIy8jYrROBI1MAzABjeJ8YS6tVArc8ytEwTnpEefYOrgF43kpmmzbnk+rqbif4A
ZpU3BEvTj90FvHwWla1nCtvX87pIrDW2oJWvDjmyIfOiXqhPTMdnYuHSnAwjYLKy
Z78yOoUutXbwTNMLzIZQdux3AliFb5z8m/g9WaouYkM4EfC6GNld0fjGQs+7ZcSD
yAcOo1GeS8JUlBuJvH36JMwOnxdY7QBW5Jor+uMrsIP5DPtq3VGK8VZidVTOQRlQ
Ee+Z3jXVZjfDrnsqxbznyzB3K/lkQBn8cfMvvpktYqYoCD6ZFX81QWBoJ4pnHg7J
RpQ799CczfhLLVNwdTVYVuRE6ykxCv6ewDC9T1ACaHRT5PT0QRjFKGBFzL7hJvML
KAcm/K8rQoV5rwyWQAqic2dYNVIqT4WERV2DIdLUQtY2/scpRlgPrx+dwaAYsRRk
JD2rr5UYzer1KuiIPD7IAr+Fz4vbpPJkhwevR39HfNIM0pXaAwQke8VIwtZXC8OL
vjfvgghDjIP03KBdXB3E2K+VGMw+0q11vJAAxK0gsYzeuvvJ+79BVef8jOeTYGWd
1+Jz45ffh4cxpwzo4qwdrD5hP2eJRH7nrU5TlGAf/iMkYWgAGZvYOSCP979KkKF7
3cGmskztbsNv3bgAJ4kGA34vA2xtaNPEsIHKlJ5uficTuhxks8jn+MpwRuAYaTnt
RJr8PtJGTGMAQkmV5mdOIMnoofikUHtCjeMXea4Id6Z76ckay0SbAPZqjc6yu5qx
j7MHMIvpHX1HBA60jMB3MacYdQjuhTR8jY6a7MLNOzHjg4Sn6xBPyZ7kpmXy+SUd
8haqIvFUOtnGdSQbnDAF5NVrgdqyeGOXyywvrE6wWHI7hU4CcwFKitSj4T2+YcEv
rEN/nOY2osFmsc82GrNBezP0C6Bh2KR40hedQJs9IFQdTE7X7fuu5ZAHsddXj0DT
AAsRsr1s2UbZb7LhJ/YVWrObPW5g5EWQgx+In96VuYE8cPC65IRnLQe2T9WlyJzB
oCrDUB9goKUDAZReOw1tabueItKtgth0Xih/GIcMQOwC7VJPhpfnlnpZ1sr+0AiY
G+bRydsmryt/4ZYpbqKRUqUZgJ8FfYLC4lzy3lSnOsAtaAJiYAzWr5FkkBZ0QItb
Yys5Gc6ggEAdJy7Vh9JvQHQmX0E0CehzF5dPN5+7crM6D4whwvuaGxh30WW+kOLg
UKMT0vidrAqq/sXOTmLZbR2qEpAOXpNufTm0HAu6lrEpH5a25JXMON8pHO8TVDJt
B62NnrGpSDCp+qmv4nxez06l9wz3IgabEQCMB8iafJcbkws9g/OhcSkB4k6p6Xa8
2s69eC4v6xmyTvlqAKJkmy6JaUSSYNO+OD7hk3ZRoF1JSJjo2dOHz8a7KmMRxwnt
cZHLFTmFSzWwRNMi6kgmZtErIWq3VnMXHwNIg/nkHfoV6hjk9ij0uMJX1ujK+OoJ
8thEq+94+8yMi2tb6whRCSmLLW4pzYj+FwxotkWj/YXw/o58IxOlSMyIpiX/u2mB
0NaJIo+W3ET/AdKy1S9sk4EtlF0QvC2o9/1k4NyzsMxM5KP1Bd3CP3t8/iilMVcq
khlmvnYcFUEU4xFEnrQs8x2tyEFkmwl+clNkIowg/qwSBiIAuYVGvz8xFV1jKWQA
1AmYpgt+kKFdX1nObjHE0AVNmAnMyPyIBbHd3yMPH4w/TQyB2vs2hysg22YnE2Bw
zxOnTftI3vAwdWY0wFEXar35u7hQMXxf5uyj5AxB6uDV/WlwYDKhjkBUGDKjjiXM
8af+Gt99BZ9PkcOxQJaVj0Eb7y7pvtj30m8b8hwOc1NrOLKJ2vKRI2cBp3R6NuZG
BfgcjsuXwXcNTapf/UEYjOxy9Y66TDoWIUOnhf5AFQbEfD2fJt9RWn8D+bUMprHQ
nig4M1ELRu4YKEug4m5frr/1lNxTsSNR0FUlokKnhIBCrFDMiNQcoZu2d8q5mETW
wVO5vlLKYeZ82wuZZqnzlYX12OInLfshvpH64Gxq3Quz6q4wYYCYz1PKtdnKwoqf
BJAt3MMNTryrCUeySUwgZSHab8ykfjw1F8zT2XyKV0py7tCzdAcFpkrH59yDmFtz
bTFL+KddJZ72FN0dODdebBb8PO3oa5oWAlXhohKuB6k3kjDgF8yMdJKQvGtVk98y
1k7Ugm8efnbZES1fSdzmi6d1EzeERjlXbS4M98x2QK9Mih23Uy/NWfigwnzwWoKb
NLDCnFslENxeEuNEUN2pNWF7JpNzE9ent74X6NB5AtB7JTqR7eeF+Cl4IFuh3BFm
tdeak2IkmE/1ZvEJ7gkaLdaaru3+7X0XLWG/qNLgyUw0tePiiYlY6w/XzL6XEvmQ
8ZMMOtQ47Csty4jhHKpSuVKPlWMiux/VjRfcIojrXtqiFefpSexDgPgP9PNiR2f6
jbQ5sbXl4cPxkkSgtPBuLzhOH0Tl4VZmVUaSIH3YnjSvO/ou15sdhHnCMxsZZWhR
In4HIBxA9bZ7VwzvYcmpEwOXCzmhA7OiChnQE5Mks0uZ61wyWiGQfpPBzCk+nrdS
zsJCNEEj9dB693JX6N7tmXVrqqCbHOm01Eunl35GslL3Wi/D1tXWydV+TDqO/6gy
h+FXosGAesrh9KH8hfI8RvuJaEL6ZnLXNiy3Ykrbl4xmozALB07gNXAVhUhTMOBz
g7ZnBxEq2zx8cz6f0oX6OYuvR1F/ogVgF09AYo/3Yy2kVadks/LVmNwi8Xz1NX1P
CybeWxZAWmbWQnr7XJMxHjbdxufbwxSdCwVg0w8fOnUA7hiTT3lOidBFu7vBqanM
1w8wGqCrhYVwQ4G8TaMWhHcdRT6bNZ/Kt4bUexs7aJJ2NGIHrdRaLDWOA4o58eS7
JfNocx5BfpUMFU3JDmuOSzFf41ULcapdWQKAB86mfkLl143+Yy6clQ27Ugv9KfjN
z9wy/xP/RcEjZ2r6HVyAz1lYrgnGpxYsmCeLQ1sGceDazPlV4GPARxC8YISbm9Bz
/8JoC2C5Ry0EOW/tQUh5TJ9amo25ednq3gfeEn4SlS+giXCj7+7JSXl/SmaEfo9e
p8DmMyiM3pTnRgPz2bomTHbJSs46/YAb2OTmyqYMVs5IkWt5WXAOu4F1mpkdFoum
/pmFaN9Q4XjKmbLW3aUXUWk9Bbxhoz5ROPWYh6u2qrlzOTp5DpXJaM3/HTdHGCmI
PuC5fV4shAGWaLy/OmVRydZPXB0Ty4qWuVmZuI4gCVblA00e04L5lVvYo893AEOv
qkdO0/1Ab0tsnb9th0omR3Hg99xkh9LYHCd3MJ/KZjOF9gjgQkR0zgDvqShtvKdJ
wecYLmtRxlF5+Wo7IypCr4mjoQ/92ILxDPAnaI2q57GAn0M0ip2JqGfFccMO76lk
BEw6ms8KElWlPZ3ONDMXiXcOpv7BDVb2Zye2iAGQahPG9yjFmOCeuOQgNNk9eisW
UR2TQXgjbufps0qstxFthybDi8Z5z9bvkGfS72WzV6o84R2+QdkQ7DvMaHwf/08F
EdhAQEt0ueuwoKDtR+aJUTQ1kiob/MBJyp07J1zV9N41dVmS9CRD/J02B5qGjyRO
xjjCZj2jQOPji72iAD+PRmaGC+BlJQCdb7nggfuYqiuiOSSvH4IrzHWI4y+QXiMg
iCQytLv4E9uHlHUv3fO5uaTA12Lzz0BB9dKFEm27Weu+ilNoYrc2nW99Pv9wjVdw
aXIRXDHUsv5IoydtJSONWmTUVH2SBbomKbmR4l/hEnzkF+na8EwzTJYekbfSYyCp
o53nNUus06YoR3K0u6DPQRqU4qaqMMD4//2ETO8Ttp+TvbhbKoTrzZHQEsH446AR
n8vKezukq1e2hNlE7bWtkZ9E9HOD4Tx4OP1FXddq8oPVObfb/uO/jAvsV/oV7Nnm
tfdO7j38KGjGOc0tPaeHFMz7gHOY9GihP260OQFedO85g4hNJla3RSFnlv+CYUw7
a6ePLZWwiahZSSKJ3XdKneXsX5PU5y2GtMzHEbceQhEsB1So0J3PJr4SI/S7N9dg
WfAdz/AtGgMiiEuig/vfzQxc9WQbcVZgpvij3d66ZcwmzrD1gCyqrCYiUdTPmUI7
ct4hxhHlb5rE5bh9l+BylduH9U2q51PR5QHkXjt10mm8w3IHhgA9O7ACZ3g/NIPh
Hk/DL0sNKkk/OcKdCVjVGLK8/T3S97TBN//jsOxxpLarVS1TllUy0GOFdKJAqdpM
iK+9Bnf6+1JhYY5pKD19QCwXV6vyUeeas2ogpvcyc38D3E/KxJ8EP0eAxP0ezodF
Xx+QjLbOjhYIae3SFnnzsI6IFjiv32l+bh+rilQ9rsIUgTOFaWnAnarJD1K019Go
eK/QE4GjIkVXnToNF3EnSv8mzl9B0Rk6N5uYTkyajOIj4Y2ZVGoDf+oEY2gCEA3T
laFon0bi69wzEffsrspmJGa1vTwhmoWK7G/OKG2oUXlVEfdqltuMNX/nfUunnjZG
cNcAhlSs9xOq6wNu1vckTe9XL46z2FiwEBrUdKyfSq9MnkMRm98te+tWqnfr72G0
aly0/TqHAAnSGcB+4erHDPX2Aseq+QSEZY9kXu0wArYgwz1RRpzI87Cd/QKm9TSW
+MQyDtUsnqW84SAma3R2/0TN5leJUmAMit5YScoEsnrfcmG0npPGIbcAbbPzPBi/
VO8xq0C10jWqCuYRxRpqgZ6LyzDR1GNY97qOsSbLZ9pVC/kGtht+i8RKoSSjcGF6
kb0W/V9Pz6yYsPUSeLQYq2oqHS8VEEImieFar40bRCzkj11N3pKRfQqYu0EIrpUN
hoFRjesnCQOUyCa1m/sOzdOabVVUib+sdqeO41Cggl81O02qcD475FaAyvgnNOft
2jux3Z7KgVVcbAfd+dSSNaGnZ3iZSKwjevB9UcujYMZjJ3rtG9k5QXAjgL5xm18D
XfxwjneinOF/2wmhLj25M3B2OYX8227oEZbdhux198zf/L3xeHmw1O3KcLY7BlTq
sRAhZMPC+kl86qC2E3JGpHpfC5hKt+2UfgwXtzWvU85NqsYJJN4vcMo8kUyWqhES
fKLLzriDr8hoyEZmSkZ4cNjtJyuDxe1uvBhAqiQT7nD6+bEqnq9d8CscnHVW6a//
toHCu9teO4WwkKkWfDHBwDSL7p2v5+Yiyd1r/cYDlLgwFNnd4Y8LO7mJVTdwFe2R
CDe8hQFVe4m7i+sNJ0Q/HTsRdkabEKiA+6sghjzQfLwjRB/Uqu2JCqeB9a1l5yQd
E2hxP6Z9Zblx3V5t/2DwPnkK3ccT/9CxrZ7nXQQh71SBUhhHLIVNJcCKXVhSaWRa
Ikd6fBNVZv2/VN9f0rMA1O+Bhj+WC8evNOJ3/6/atC9Md8Ce+wOIXYLwG+XWL9sG
GV3nEMdFcoMMSIS5OBofN806UUtiJkVIRQNzeCNVyO22aQk4rx565qt2Y8fw60yx
t3IwgeHFwy5r1lco14Aggjo7E0OxsveuKnqC0mAlkNTx6hYtzbrLw7luoiRLq220
ure6miyNodLyv2eDcasAHbpxi0kl5EAuU5TlmjwWBjb8ii4TOexfqD2MjgMVERur
HjuGRjI8q+HgORBuK5h8LPfrujXA7TCtMeh4l1aIStT8bshZlTwtn4AwS+rC3wOR
nANIgR8JbmBiSyP1eSCYL3jDHZRqknkbCnGUgCDYulcXI92g0oehdV1momNxVOSz
720DsgLhJqkrIL/q03MY2AWj+4XMqOSaGLTDNSisKzAUgwqNx4RcIkV9CPw4BbkP
oPi0jG11ygXyrQmuLEl82WywGhEXFitD83pP1V9HMBeei9N4X+BAB6M1JOUc7/rg
KN1tLb+05fLihUFFwf5/1GUz1dtcOTyh/Vs0hhGWw6fma8jdxcdZoteberoElxnR
6q3t+OTqCQnqhzM3Am/A+S105X7hDOzwuSJ41umMZFjR0/Jp2tPlUy9yOxDox13d
O85fnlMRrkkq34+jQh7kxhMbXdofvgknWqiU0qdrNkJZBU4Hwir2y6Le9MsRCovk
RZqfxrI0kVVOJZcc0SOEb0ov/KImPTbT1L5wIdCLmRqiSeYlZIN2JcKeVJw/MUEe
u6h8YMey3Cp4drd0at6+ksOxzITqSnJy+Ib5BTrLyIYcCYTkX3HqjJl7cFrvCqLA
vZBPzYTg2I/zJqUThXXQ+SAhWCd9gGFZmKA5szxWOQYbprfiSSN1hyRRQfZSn9I9
z5I1DOTCoLBD8NAlia/zT7cC0NlB1Ve1dEdLuG4c9WIE4V+sFEbj63pDp6AEty8c
kE/sQy3vIoGFb/7U5b3N4ocJifTNMovRNLg3szMakJWAQJFBubiRkITiYd/wGxXT
lewx/G7KUC9xCdG8NM6JkmIFKWxVVLzGwGhFueu4gdV7/NidBSvTQXfbpCaNYVHF
dwiSQz8BzxPCe6lIehWZaNqQz+y/xhpeZ7axjWbw3UC736QoVeeg7uQdMYqPMvBN
eXMuNTXYAi1XUJ7COG0XuFZ1/IvfBbxxu3ONgDgMTbizHZ/+2e4BgikEdb1htbtF
01HZNpVhf2n2FCFUZ/39xfV7+hv3kjKYKSFhFgAWt8yV9uOh71wvd5/RqnjhP15F
jMRxT1zJMRmMDoNIJfn27wuL++FldT8Nni0nTp4Cwxlln0aO7XCZTM1AolB3Hdhm
09oXEKoqXHiNb8RUOPi/0Eu8/tdViAup+wF749csOOOECQzSwC9JnKHRaxfWt55R
FchwXL+zj0HHoJgoeqZBtrJRQfhqIqM6wbgj/gEFG7mS84OOGJKcTP/QIpMvyQC4
F+fW+RnV+b2VHJLwgl62KcJHEzWBraaDgHpUf2se1r3eVvWesY0vRznQgBPHFC1J
s9Q1dRX5yfJs05iw7DtScNuXU3fam7/Xes7JGJE0hUT0kI/Npu/ejRJ64f4K5hlJ
VESc8UFojhgh4TegHDrunFRfxuor6vOvwN5myWSApAgITfmwNp46StxfAVIyXwdI
gzT0fhgWGzpofYjMLg3i5KAbgTic/on9e7FDM1xQXvLdxoORRiSG8f9wVegqe4Ui
jworWud6t8UmjyL5WYgBKSquNN/mdHmdUl6KiSyILyQjZ6hbRyRTrrMPOaqipgpP
ovhUNf2JgwAQMhT0uapjmwb8EvsS1flEkZm16cNpqtGCFF7fEx0+paq1u2cPejSs
vTu100eIsQQmZkWFR0YRMz+v4Rt1IMoTldWZpETXBQ7iJC/b882tAVGG0mwXINCt
oky5rv08lFaDtuo0vrXXVLKAUfplDJaEsZy/8g05HZ65AHKE2r8kaLpV6aXcgV+l
UANArYeF2/pqSfDpKzVyfSjhorKFZVn8Z6awHQCr2hVZWNztCfX+np2m3FfD9ipX
kLSVaT7TCjxx7mWKUBSXjOg1GM0Kh5FPEOtdux31a981+7qpG6Of8yosNwESWEZV
Zmp5mRVuYdPcYxS+kaXr1Rc/iGHqS8dpJYuNbaMgv4sZks7tMK/s0sPMUABsQ0e6
tq5DJak4dxydWaE8llyLCHWje312mjk8+r0Dnl27Rlg6tSbxDsbfFCdbIyZFGE3j
ncdXFboshPKN7kJjpF3RqhLkRCAMeP7E6LwsVc/sXKvzAcDmkQhFdnbORN2y8C8E
R4Ddhs/KqlJrRWp6UenRzRWNbo6aCWRj4qCJFA2d3GTeyP5gcL4MY66lT5XGtFMQ
JxuystgRcIw+n9X56bqGf4cFIMHPQVENHnzSvOVjSiKgxCh6srf5IZiF5pUJJUwH
Fbaa6F6w6X1Rkn7bXNnE6gqxBCViqtphgXuk0nu5vLhKCsy7NkpBLDpUA5Oj75az
IF+nLkdhnIGvA9Q4WO5WcTWHt8z+vIXacAp29TfV+pLmm7AO2WFzqo3cbzzialwl
66pXyi0lX24SWDPmogTJvfljAK8DbQfAMNweCIB8Ti5yHwyYxOJq0gcJ1pqqhDot
w9Y8+2bWdQmsyTz4V2SxhGaAKyCOER/1HmkdFhr8WU/jAEoQO/00eV6ZUEd0MISU
hyrGUofC0uCkIv3kUf9ql+Avxlao/qyI7m/0jAR6DhDyVmyeKxBgvmhLQcySAL4s
8cbNuzjKj0lGqVP4xoPErSdLxjYdcfm1umPMYdKm2xRt1Oxc66sRsihRLdJ4nGbS
UwZ6TPOxRC3JVrH9ISKvFf6lX5G4ugVLFfyPBXToS0pySP2wmwuiCp14f/n5+rBf
e2jsXBl/HRhZxUR418mspmRTr2Gciz7zXHZnbv9KXB/MesdkgCvgqtHpazExuxJ7
MFHeCqmvGf7o9VVlXN4rtNgDSzXNOX4spjk3komGO27C3kK1h6FiDaWJUOlyMmh3
A/EDj4WwxDOZ/HVgiG0cOb70RaNITMGV5n+Y81O6bLHqXQKrDG8AT8C0dBy2yMDm
dbSoED7553VMiEraXIpCJ1tdWRAdqmpV6bZxx0m2YEhYQusObhNtUpg/D9OhYe42
AV0xR1Gq8yYn00Emp/tn7KjuUGpZjmCIYHI8gegBbsTqklwPV9igqF7Wno6TMBpz
AbZK3x1yZfWPaWMKLQm5E5mun0cwYfOH2DyfKazwbQCd78QA5VEczK1fe8yDZ7Lh
J/7+FyjgrdMaWeItwxAgjZZj9NjwHTNyrYmSyYMjc6wgPY8j3iZcJAI33OG1HyxN
eEOINpPG2lHWI4F+/QWlTIze3JH/lhV5nJD1EMay2J/hXvye/VfDliKzkq52pxb0
kPBxqWw2+Sc2USJZfTwXN7i/x+2J8hmW1AKx27qvxfQX5Hvd7wDpzOomTlocUH30
f3ofspE39RYmW+t+zdLrpW7W3SOeIDO531ANd4vyX2f65nYVxn6knit4yoaIlYvT
D3XRm0PVNh/5gM6AFMR5JZEPZJaONac+9p3TDiASZRNeBlOncJ6ZeJhc/2fzuhLe
IIcso8EDPR0qhgiHsyf5kA7jI5Fpu7qTV+NC8sDl7WAm9FFXVD7nHXO+6UEoUqNR
7mEXphipb4gCUFz4ITvpV0Q0thgSP9u0cUba+mi6tB6H5GkApb6dCfgdX++HZW1z
fJCqpoijSQqnWbzIaJhIV3o1PKdcn+nKpPjGZH50RJo+cTIX2tgSHPW8xmyzqkoL
FY143kMET/+F7eDANt1LHqfe1TEfRZ/r38f+q5b9Hyag92NlbKDAWnynZn/NOYCh
7PsNMRcmWAtxTx+dni7YxFLbVEqfAuDCK+dNuuiwveG66wRJ5qTutel3cWTefkQN
miHDFAO920NrDGI8PWDDi1g1St90oyex6NVZj1kJGrOzSyiV06xsodjzqjOv5za1
QNOCgPe3w0Xq9hKntd5rk9N31eozqO0pf4EMKg/jmiJn0MBIjkKrlCNODoZl9yrQ
ORRzkFjMiVHT+KGO+e7zmfrCsh1P/CLKzKaFNB8jR7G90gAPdGNktdizejQ8HH9f
fdZJ1OfEqiZrHy4VQAl7fbQMj0Vf7I/RUUBTfdAyTZZHdg3k/6KQ738FVzjZAluB
9+hhPYK7/j9079aHQhDkPdpVNefCjEomvUGYSC/h1Oe5vvYKHDu+tkvxeRZOVrGC
B40zIQWszMbBDgMO6jEqH6AbfGgIiQOmQZWiNqA7qCeodl1X6BdLaErD4bX82IXN
dui15WiWtalO9yqNtb4HIK3mIc4Fl0dQYDRR+c6RvbUGw3o6BRei8R/3dF3OMNlq
DBmP8DxK1LKv2ShTrvZIajDOoj8beGNU6pH6eBW5+3KjMQZ5EClkHdIVYq133yNZ
QmetJPBvoZvYmtbAx8hwZ/a3mN4DDes+nKea9BdN48BNY6GK8ZOSjnsAbRnyvc1V
wz2RZmew1rdbaC28mEzfhVF8zMVnnCzM7GeWEaCWCnIsBHEqbbgixXGzjC7DD1jN
3BxdvUYLUpCN5ZDCEwQ5DoDhCOJIpvPzGm0J7on4LozcqJjzDAD7cjActjwVd+1Z
bp8uVd0JAt0ATHoCM9A3TVBtL7z4ir0vnTUbjitujRBa+mFMOmwiELnqyoab3AWp
h1hJFo0tliR+LttDr6XvqdnpwBdwWGewKBgiUgZDPxYQFV5EYU6Z7E9713UqvhG8
GRtI0iN3+01nXaKXEEcAnS1hX/TYWF0V+zFiw1yWVtX5/C0ETbudbyv13MjkdaNO
gUcDZCk2hZkljyHvlQ1Chi+ZUMak9ijJLT9ju4wciK/7sYGI0aVMdmhNRzNBHiGN
OVVoDQMRQ5MKiBPFMPtk4v25ZMS7Ihjb9Q//r/L/3KtAYm9b5t4UAjOdAT17IlkU
moFC46eFfQLQxGYUvRO+JmMzkUXZ0Rgn3imw1B/Y4jyDrxzpfuXxb7wusJSp/GkV
T9gol5ybpTtkwCaFastbuHYHs+Q3dt4dUAsJjqETC3WyAHAPR7JoVe/XAPYOUeo2
4puLcWQt2tzImPmrG5/kyw+pTzpIwyEJeGxja2s4JpyTnsjcJfQN6iNY8nx4ivlE
LoRO+tgaPlVkOF8ItrtoVq3fBGb0Eo1isWPJH0OfK9g2sWhRp75XVKEN6EpT6bh2
bTQveE69PnLFOMx9PoX0ggk6InorWB0lCb/AicECdybGxE/QSIoxbgrT/dpry5rC
7J8TuOYRz4B543dEuHD6XF7F5TEEuddMsPpWlp/3E/Zhsiie33LkP1KawklXNQ6S
FrB6GVcJjqyNLTFj3jN3ykgbZYQRkbrc17A+C6TkszX1KTIW0xd/f7GkNvR7UlaZ
Gf5m0MYQphCF5KCMzyn5LtS/GwRWN9rFGKkyzGrJzy3gPc2b8MMz3L1vFfs88vdb
aYuuuFSDWY5qoJkUHLgYOwRi72UkQ6y50BtCqjFS8VO4Vf3EcRtA/3cb1ISXR/gi
EZq/k1P9ZJFj2IdJmzg/CMGSFEhcIe0fJRkJx+3DqFruMnXD2NwM+7Tkw5GDUxPO
u5vTkXo/1RdVZBMC676VxzI+y4ha4fCtbUr96UjYimptkW13PvGM/VThHboEWiIA
FTTnBFMB5oS3nE3icnymsOvKQJW+c0A5YIt3PlYzapPYR248osjZa7tgX6JZ2FZK
VzAchnHr4ezy8gFImwFF8/26x0VmE/DhVxeek3c/LNQ8Zm3WVUBNJTYACpsAPZaS
VJ4sK8+DjkHT4/3oIoyVfHa5q9bboY15nRoCgM0MJ520y5lO90wTF/6wE2w+PRZ1
I/qpISVKq62rmaD4oGKIwS456N36ZBZvjRQlCfrFEEJCbyY3jqA6up6a2Wh6hrMf
52j5giQDYDMC9lKFg+vF0+m5lNFFPQlwkvHL36oMiN+o7qC0HIrYXYiDPfOIXFeE
L3O4p530ohLYXGwGMAg5ep0BIh0dJPdYKLRYtJ//WN4zC9WE1GCLAGVEFZ5+uZpy
d4ak93t94Uvx3LsNuTY1QY7101oYvXrnVVXxKLwZXQjuvnFlGj1Yxs9k9osj8n2P
JJLlJHhfRiO5rCblhGXTRLR62u1vy3k4/v3tsq5GWW78/zaMXaBPm1FiQJ7B7XOd
aPN2SFBmDKGfYB1Qylx2Tm2/+d3W80DXOV9CNujIoo1ejmGoXfraoCJAPKsr7+if
Y4M5y/JDT3n+f7yijcpAEukslNpvNrUay7EihrWIf2kNXSxAAM85sOtYWRsBRO/r
zAcGcundlejELsLBJ92Z01BHdcQtATNRlxqSqUhzlmo+ygiAqOdUaaBP3nCxWFhg
tv2qgOQ7qH2PMm88yiTOcQZEz3rahRhM91JsVcetv8y6iBJYvucKLnFX5903haYU
XI3GvDU3X+6Kn1ePCwZPmd/JXveGW96I+Y2R9ISFpiBZkoie1KZZM6XewLo8g5Gb
vSE2bM44ifeMCYhgYLy/EUMitsHb5Snyeb8EX6ZolxRqHg0/OcA8ou2HVdvPPWAI
wlBNAzF/fbhqNW3RA9UQ2ZVKTItj8tc8wp7ivgEDVOzrYAg0r3Ykkm5uKyu9H++j
LctNEXw3UvbijQQa/kRlGz2jrbpMB0t7dzr8inXZlY7P7MtQyn1QcorMrxVRj8Lu
6/9BfYYlmnEjWkRteMWG9j3KkKfIZm8UEo5Jl4e2UJ7SiFajHnUrkT8q59Chl+Ja
52+viZIsHcuFI3PQA3MTkWWvKMpgljfgkrgKRjMWjaPxR9QIKld2v1KPi1Y7WRJ4
9qPmzUr0GvC91ECKCBM3g8a9FZX9y8/I2f+1o4zquRXQxmg4I6V1uCbWGGlf74M9
AH8uRqOik/SmRv5K0sXpoyMxuqOT8Q2+6faZOH5EfoKjUfe3s28w2zgpVhJMgCPS
2nkG5YFQF2OVVAxTslDiW5AfezXQ4POFCtCpUotWkFKbf/1NYoS5fXIuTVlFG/ut
/8zm2FVSPMQ7K93vR5J3of7aR5caK6Tn37BMMEKAjw/VID8pZKQE6DqRum8YxH1j
fuD5PUKlQ5+tau5lQDz486kBGGP/4lXOovo4iCgGJGH3CQvsLFwdVJ8XUiMd7pLh
Mb2S7+sehP9XN/6mRkbE3XXus1nWE5ZJv5F1rNruRAaeTCe02+1qaH3QFEcRwsNc
+DfHgeX3qK/KozxhJq1zknN1TEpy+9VatFzOgyVSGuEEKKzsgYIINUV6+maxs9KH
WX9n/lv2XBAAsyoJEgBVT6GCgtVfI44b9r7Tkj/BUJnjpTKSTm95qa/MMGMeJV+0
RAKcjhWq/wDDKaJqtojd5z/sVUZr5vL+cZAZKblws3Km8OLveo9E7uDnLfBQAGCZ
782sBptT6ima8qzPU6u2zMuv+G8q5jC6NJ99CzbDSTm6qyPvyTO4g41f1UUwzZPn
xgrpLZ8WwQq2P9H7+OsrL7N6Q3z9Fw96R5DTFIOe/4XptRXMtuj9nvr78BvoJ/jm
M0BwjjK/TJjcAsnbCw9O2BuIuWWe72/HBFipioUE8K/QtRnw5n0BuvzWAp/vGnCH
+OXN9+lCro0C/XklFzMqnQrDm2hTXnlb6sNygj9KrEK0MDRSn2+dxrOzVhbyqm6Z
nlJ44mckmgs2mAYkK6kBrlbUDjRqrAcDsBzREdY9bvbb+rSqQ0uY67kvgVBUYPO8
U8XieZmFldYSG5qDmTo5px32oi4ySi3C3yARXuTZcMpy7hE3nc6oOVIieTyk431K
7sDWnrzKxhutdEnRuNlLePGsTJlzVu1RQ+CX9dJSvvNCMOGqXeq8Eu3OOvlNJie1
HuIJj2f20wnx6FJB5DhyvluallhfyHUoqzBh+5JRnJPFU+W2GpDTIEj21KkE+X6t
sUJJEmEhBikJNRMF1WQI9UrgOExHe1v/qBtW0Wn2VAgUdf0Rk7fvQddfLceoOoGL
jafTDVaQh8sGJ+oDPfMdIfnfRDfbdmjPFxCXHOWvWxjo6PDYtYmatI1J6mhAJJXe
sClLm/2ODEV/kTdZOq+5VmCe+9dgjdjzvJnOhwfIOHv3BFOzJAam1ISXwXnLfZOA
0k5bgaDF4CCvR7reRxl12vgMPeAPjXtZbug7s3GChJqhI6KqX+5JwXWnJTOlLxAo
F5As2yQ6EVLN/HuHpZo8caSzsHyWQXHcIC79B7Lb/gUHlJsFnJgKtWrM1WO8LajL
379orzP0kVlZvoSo5t89FMDuft53KM20C22PxNvA43kEBKqQt//2cpqMwKy2VixH
6qeUSYceDYoYeVgmwBX0GBLhdFLbJmM0YqDsESul7N3zGY+jw4j+QVAzdNMQkq54
wAl6OuXIENCs6ohNUGdqbD866J6+OvkHdrHszUDzD0IqfdxmnheyuwcB/OOoHLcU
FGXG0HlJQDdya5pdwrSdrEiacVHfacqTPBNxhf5ha0IAgFPPBrK9R0oW1fyWfEEm
8+FnyOMQFTeOfroPZxJsXNphRRYG50Sym2OKpj2YqhNH332eCCvh0zCqvWkrdxdg
cuckCsfYtQfp9z27riHHj3XWK80iCOr1qrJLyVPOHPOHLQ1cAVYPKKXnNcFDtJ0m
xiURWagmfVysdHTQKAcAMxmLRvRJnrtQplBFUt/r7GqdYf4Jsry5G8orNeWRViW6
cVZGBXwSC0ANHwPzSDL/b9WzBXpOz9hnXut+NMkB5IXPQnfOzYwVoSalsfEU7vG0
jojHsZ6vbLD8OjiM7hxud30cs4eJqujClplY22q+viv84vyRWmVRkSw23zvJRxih
po5n7pdRVh8BSm4Jntux6Tj2slN4jCwEZGJbf9B1w+3i73OgK0Z1a6K2hGGQBdM9
u6yMIyaFf6zmLmpJYg9v+TsjMcdkz3rrWsmyv35zD/YYkpIWBYa4ICRhoPA86QrG
B1+D7bj3KmjwE+4ZaxAvAu3riyAxC3MgW8M4SnoyewPnEktA6QZOrlo7K9T5RdUn
Y2y0OcHRWEbhlTBcFDfW5tGpLFfR852zsSNme/W7BMUNr1ohqzkHBBhs6JDByCcE
THA9+W1Vmmu6acKq2S9B3qS3jzW7W6KFUsSJMLlz0b0f02dX/M177GqUbnhuuHuN
jc2MdR49gO0a+CmVsQxSwMK342IiGxqEB8+RDQgNL32bWFkMfDbYYib/S1UNUoFN
UIl8asX5xeGsj8Ey7OhWvbKzYBnJZmrtBZ4EUZx5uAAld7AfcAVOwo79GcwhLGEs
ECjZhHGgRERd0DX9VXUodtrVpS29d17CRDrPc3c6MO5EgtwzQZDlVMlt6DAAMxYm
qjshUPL7h2trwEw3xUgU+1wq74I8uJvqezl8q9oWAojZaZz7RbxMnB98Z1PcuWmK
GCxdNPmjCh6K+fKNRTeZJaBMFNVlsNy9pxzADWSTTNmHphsZSVLP64IFE3rkJbq/
vJxDqEe2A6hQmhC7EUOCFE/roogdPo1auTHACb1fR9w9Bl96YlsYHKUprS1jRzLX
YPI9vHyWB9hgPHXT5fa2n8dvw7p5YHMEFrjfeOxU/jhYvISptmp6Fl6WhGG98fgH
db8O+8fk10uLEKCDlWVM4UZeycoDQgyn513DAKW4q5Y5aLpeD58J5dVHI0ItPPPI
J08hzTv8sImVY0jOyP7y7mHWbLrL1BW/bgfr4BZrykQ/pXM/8OmuZqfxmo/tduqD
QVn9WTROopXq1Ci04JsoSogDjWssjkt/xlA9x58GUTXhBUe6omVtuNMlrGQGe/M+
uoHKkHgAUAUOxay1StanvxUJQCmG3a0FFGQzmUa5sbHLi70i8NOX9BdGagmOL28B
A2fBfLOIJzTWSnxnwM5xJ+Nln+fmD9/QzCLLV/QnDdMZgK0ag8Edq13uSToR/p9d
dzFmZTkUUcv1/sVXfZ4femav+cSctzf3WBXk7H3yeGRVbxqu0qJQtG6zuahs/zjz
kbXT1UtEP4KeK2g7dntlb9RGmNLckNs8iqM5okdQ38yDuCgZsQM/xrukmGRPemhI
4csxK9GqxiIS1NGJIT6sIgvn0ZmAmlpc85dEfsJLGYFfRSpQEpWwfJrw7FNK9JuT
2AZm+hxOJUu5CKKD1do8lRcmRpEM649zME5y6Nwz963P4YVctHS4UIGcF//dNktF
csZeObRcAPyD8a2WyiPcUsbT9u5MiV7GqohtL5q4jY/RlcrHHnHTQuhQM/19HhoZ
LXvlwEeDVXK6pEEDAHHLbagSP4qxqv07801IHBpO3Qh/rQdhH3ZD8MaQYMDqa1DP
qkEWB+PjJW7v87LPMvHVzDiy4W2g1JYrdgyst2GH8YpzNSUy61hpUxWA1J7xFFbq
WvVBN7lrFlR2am1Kg1s2btKX23HnvQAR/W7BzwO7Fwk213k881UiHDgbtkOF24G8
K3MWwxTT7biAFUAd3OBKRlKF+TzjPf2MpGK/xcFFeEBcOqbySEIna7pGnNKPWgws
DDtPfxCeVtpVGFNGourTxn7PGt1y0wV1DacBmN9O0bRgP7NaX03Oc+FH4daKDdG4
zbu3YXwSQL3jl5ooEkNl3KUFAg4+lPrqBcIYzH7k1ivefCS6tZ0iFW+tduLwSRm3
YkDpomGT8NnoZHz0qRajAYORNbFydvPzyvcE04ZlsrhMl6EJLDxHxzyh95W3jVMT
HzpF4XE+gVOf79RP4nOJJ2Kv5SgzKnkmuBFHM3wSbT2rgvWI14kaTxVKrVG2Ki4R
4bgNjUrAK87CNurg5AF0BERTnTKNM3NdsSRekzK2wIva+NB2UaAU+SovbI3jQvX+
O3j7JOGS0WtjFZoJfvVLBUpxbSPvtzYHNh5ogk+eyRaGG2b5eWu+C5A/wNYVogWY
eehB3m8cPNVn5QO3Mya4yKDrWNN2Px7CfjXZU4SgbgTuUOEY1bHFMFklKX31V+5i
OSyaBQrfhUmeUzxMnqjLrugC8sJjA2gkO8XG4VqsjUMq3sKmv7Zmz7wI6f0zBEPN
/PyeHP3QAwfufs7Befv0EMsYUv+15aIGLtsGWMPHYtiTbTwqk9Cjth0GmPiIDKpk
ABQYdoGK0B16UnozMtiz2j/WS2FaQEHMhvVa6NA3v+wRKpZz3F7CX+RxvZy+kGSc
kpRt2nSUF4mFocavlehBrtDdgGhnWykR121MTGEK9zUHn4YR8AtqWOZzAdYC25RR
YawrAu59Fj4mFrLUoSUYZ9UlGjGzyvP13uNoQqoy1ZAyG+E9vT2BISBSJ4WbnFur
5aCzmr7pjzxgc5SCs2lahwh0Ua+w9laJNN8MT4fCmtgTOdqPfBAxgL/ummBP/1WM
Zg85muUASbkR0JMTygQPWAlsTBPjUpKiWQthLRixvjHEgZWo1GXowERp78dr6sYq
FEbO4/aBzj0iTiKunAxEVv1at5FZtxd0Yh3axQpUEAf7eZ72qqzt/x1G5R9E+rC7
5TZqDXpr3qVf2JYTxKvX5risVbJxaIFIHCX59lmYku0g6S7pYpyrkq7Wi1i+DY+M
gxJjeqLE1vcs/IV+CCfQc50PT5VG8ccpSVn/z4PJjM//85/ZKm27AZAoM9iPr1UV
n4b5BMOYit3Qt56RYS3fMWySAWHt9kkLKiQMeB0xnaVwIodWlx4dExMDq0gS0GML
XtyHpgwwF2QqqXjJfbyxQ6Jt2eCinX2oFlZv2dSmkiYIkqlTaGSf42RqHLOhJJq+
nKqnPR5FY9lmvZE1D+IIyWtn+rdXjYTzQMlAk40gDB9NBmRFy/4jwrz8mkwjhaPe
/sxrXE3lqOM8pee8YspMd5+7ZgW+VY45BXmbUsgwZcLGdkXf2Btu+6B/QvguV/sn
5TurGHjvAU8gPFlzSueyFHpBHdAntxCbh1Gqv1GOpZTbkInGSqP64CWl6XgNoISg
IBVYAnrWcsBxzZSkBZkGcYgt8lcYwZTtMxrxZPZJSTir3hM1dClBoGXK7+N2jWk8
DBwEDAIracjUgOzLvL5mG2wPP7pLDMRFQpJANpTWw3niHgloA6kmQbKf7dckx/1j
2tl0b2anhzpQb7Evzd0oeN7352hMg+yVhtQ9cJR9Ae/LTxA41Ka5HeDye1ezEsLW
4pxgPotvDXqoD2wWb8pluiSuFziOoNuGNfRkIlFaxMdn4hmALxVjA46Jv5KPxAFJ
GSarQhz0cxKiUrXpVVga+3GChuzsVfUz/7zMgn3OrX6zUBELlXKnvMQJ6p9pttp7
Zf0VJXK0yAezi7tGbKOtp6VhJ6i8mfcj3P8aSHyDLxNgZL0XOAYokhgZpurheo7E
ON23bIJ8rxd1myzasthFbP2uMN94H8k5APci1phhwuYeBBCNUvG+d36d8bkph8Ul
ep3cO/MJfXAkzZXXF1wdS6ysvkK23sOdnq6CXEP4HQwgtn7jpThkpUwXMpgw2a/U
fxluspQ0YX61YvnWbFfJFWs22soUulP6NL+sYe+8pLp5snB0j7rxdNf1qziUafBp
6uKW8K0MKGya59U3bMrRdL8h5EtE0OaDID9H/MZm7wdYXt4eouSteH58pii7kGZh
C72iNuEd+ZduJ4R3ut5A3aFTCdGcSRTzp2ILhYgGv4DlySXhLRQXufBVUxbSYdsT
P7y9KTRMUijdVdt1oO1Z2d3JKNoe6PXLvBZkVLlOR75CGqKQrgXa+6lc0UxdLgKA
51k0leC39xepWyTiiAuBEtzrDBL/KsuNRP0ITG6hoR1KWssrFjSDbIl+quPM8WLn
Ri36j6mcasxo3JMszGwRLyFYmhUaIteC3bzMThNTpLQQgUuQo+wFzGupeGGtBfpJ
493CdTNLoG9rfOL0ZekYSmHt3t6kI47Ng5yHQgNfXN4jSwxr07IPfqboyCOUccUF
RcYAO4qGCulRNBrFPnABnsYQrQyBDQaqrj4wPrOV2b9hU/07UJIePhiGxgBesR1P
Vyxu1fKfXqYvHus/hZ5I9Kc00GnQuZ9NRRqsnzh3CpoaMh8epy569l24DPEwt/DE
ckrDPygKwSfBhNUkeY55MBV0UJXtCs9hTOILHjpwp/Q3nKaxpdH7ePyPghV4UN15
T7ZgTVxgq1/U8Qt7XvPSdYV4Phxc9Jq+ARDd42mPxhb2yLX9rntWym/sJUNCh2YV
nhLx643BC/8oZ+pG55lCJ5Ks86oEUKwjys0GP7XKIb7stVH9rl01QZrZe54oaySZ
AhE/EXK1JHsXp4jAOVALdmPHw2hCM3mnbHoPD7ZfScHbr9NEeS0iQDo1VM7Js2tc
zwm6N2EC3h9jOL4/vklraBt+lz6Wj2jru9izbZ7lpCNf5pR5yTcF3NSvLrbKmsg2
B3J6YZh/EIv9z7UJS2YCfhn4XylCPyPmrMnQozoYxIkiyBcOlnW7PccOCcE60IM4
Hj5ugmHR0nLeWjEZfqAeRdHFjVdPbcKyeMAwurTbzJy6OLVUXsYiNNs4qDxM82L3
tgNHeq7SibdtRYgk4AtbyYdGw/9vM1fuJVmg8FxbtGI2C4ng/x073e3vkxK8kG+I
s6Z3bxF4NHizUVeax1GfVazBQMIXosnd5zJfiF/IkO8sT9E+2CKd5EUIhjg1MQ7F
/swOpNlAehd8WJ5JjagS1vTGCG+fRzzz/XEVXXdbPuaSMBFz1mXIjJJbPBYOqNRA
jDN3PDwNtZVAGZ7KYiKBhDDelxYhhnwCbeDEG8e8A8DtEeuvdj4R5RO2zPnH7/Hv
waM6c+fJNg7U9Nd2KpNG0VHilhXDXHL1p8/fogFjsa5rFV37NBbnp3YXVucbg57x
YCwVIJ4unIRQTEBHEOuYe/KEvGsO4jIjEvl9kYIlSm8tJZDLlKnD9MwU5MJel9/H
doxmNZuwLInFeOkTZxQSWAQp6UaueRJBK8owvWK+/IzZyxzSRzyvOdb+WniVwIm2
4/oDJsLePa0KRcwDL4PbDccxBSb1s6njYMdc/iTmkATPNVmvG0eKK5uCVVteChDI
zQ7xb9XUpGdzea9usXXDQFYWBk7e6kTrRA3scC+PTYEQdvnk/+qIdDrSstM0gzMi
4Nen1aSoLWd6zdy5PIE/6/2irWeoZXaM9vXyFwcHRAwup4Ical/x69/0Xzp91s88
cXw8Wtw9Tu3WqJ5JrvgTKR3fGS/EnDWwEy0jd+PiqDNYT92PZXBpnQIIwNMU2J/G
fYgqKkcB5GTJOZb2z3JC+VmRvEmDgHCxaGqb+eNxKRu3RkP8KSZMQToMmgccMrLD
hr3uDyJ4x9tcElu3f0VCr48gZIutE33vatE37icV0JMNF2kNeZ8DflVOpQHdf2aK
VAVaKSwMEuB/9Pt9McmVRvPhQXua3EeCGA97CkSTcPbRqpQ9GqxWpmVdg64YOy3+
ywYviDiits/Vnghg2M7GYcP+to0WvxcNPKnE17DOBHCHtBqd6tDeee6NwQg8OQqe
aEAsBrmMXJiYJk4Wi8fZ/H/xbVeim83QKlRWAEyISYwjdlx+Ie9urVEqfsJv35iI
MlGUMQZfuCHLBX/Lz2OhpWvWL9bAUqCH5Pxf1t//xWOVGOzqnUjRF+3RruI0kDQi
PJS2eLfhcaAWjIWtAnd/Bvu5NW/8yBxY2z+xREPTyC0IJmJJJzUSPxm1VZz81lpm
+6bEOpkNWarPPAQoIypzsqvnWb8yfK/o+Kfa756SKqi1zQMI5u6Air0eNF0ZkyIW
KqBjPVNskcgRzp0N0sjLIjzCoer1q3oVa8qPlU8BNt6rkLyjN3RCWnjveL8Mcb5q
4jWCBaXNEzApVnauMPluat3hHuJMx35phrl1KDM2QV2A4XcvK94nwcfGQAXMI8B5
IX09/5faC58iIORN8CWAdeUxNisfb9BTxK0y2AfLeuvk97su2iWJDsvU4TyUvM1x
kUYIUhCQmZZwHYSG5aAbFScPXfuJUqPfcRQqmwIgqp3ICuBdTCajfl3Voapn0dzz
og6a/RiMTVxzj9X5OIAjvztnE5rP5hDRnqd5hGZBkvbCKdtudzNA+vXOS5kAu3Zj
inIzVj9DhBfBLvY0mELcypaZOjVgpxZwXslUkFkJN2I+2sYQhedJ8xSim0/z/YsK
FB8v0eRVXBvBR1sq0HlR6J0OWbZO9BJFir2NcS5wGv39GHW/ItT1pEDFe59LAF+r
HQgwsOpjDOFSDiUJVWRkQzO5D5W13nMdDZi9s62WnFm+LsnxYloEV4hRulg/1AFO
RL6INcs0yCfwFAAqJcmXWPJ1UBXgUVhLpgay9nizPI3a6+EJQadzCiEnVC9Lj1Wp
1Sjnr9Y1cNK5ARXBlFyqXz4CEm1FsF6x9zLldQoHvUU3G+3OoHk+ElAy0wANnrZ1
8IIIXAtB1Uonm1GfavTWS6oHeCklshl9saeYpDH4egVWohKoZirLVzWYalimsCIA
v2xHRvPZnfMRBLunNPoonz05BW8Mr4ey1t7xQ2v2fCikopBpX0kTirJTsG5GsnMo
HIgUvzhUUW5CVucs1mRljl63zLK51ZfxUkQ6tyCZY0oqOodSC2JB/WVEquJcskYX
d1BzIWsqyM9oDaU3isM+bpILog/hd2nSSkBwUwkKBot+NUmRVM6L74DgbMrI07I8
m5+fsWANtmseDiXJnUhktmUle2FeWklcmoGummliV3G8NYHqZzGZYg0othH7vk8f
fjakXj95QI+XD0UBgGWn55YICz6cQUO173a+rYZDnBbRd6TlpVgEr+ciNprF6mOc
sw6GddGYtjUnkJJ9ZvoBPHUa+GM6PzXrM6+8Rw/ekfp+XlP4bichqN4FDJ0aKeTe
6cs3u78ydXhHkyVBtTpywgU/nfOhp8PUScdDNL08frqALvV/F0DEQOlaD0Vo5agJ
MrlqVwODo4x550MEHe9kUkK7o38fCGjUTTHqoR/VJFFlaNEwM5aLpOu3A7GTu9wB
nrNM8Gplkz3pljw1NnjQxFSXVhwSvb7eSBEmro5wZ6SDqAEVpTR2dYvyJ6K6pF09
yxgsy8bfVNJZsoUMr8muUsGhIOF5uKPuOXIUYKwNCV8OzXym9sKF2CjQrD9rfISa
vVe0SRG8PaTa8FYKYzr809QkdOfPPY5YDxRRFlzwidwHMtjWK8PO8mRiBGsyMkYE
bPAi3msV6/i+CbyHPnEV0+imJzruz+QjvO+ByanQbQQtl3UE/q5eUq0oieIy1TUM
O40g50FRvjzXbyVha2tyW4Q5TUX8xMiDf3a4HCaihD9gBkZyeCa9046xrA6C2t8d
f2nd1hjwYuBY6odCTRKjt0l+LMIpFvwV6ORD/DG/htsE9qQWbILxgPYqIbSbucZy
/4dkq94PCFtmNO6uvVz9jVjytiuVvDtdfOpomJgBV2qe8cqJJrOznbhyn+Yuuksp
g8+UjwABThhH3k+CQabYhoUovQf7KF/vHs/pdZ60d4x0cNV5lLM1lhf9aiz2JddP
Z4cLdXrDbeMk7zLmlp+FOaD7QC0+rcw14nr+by+5+/ml8EqWJmYqPVjFKWyL1tZ9
f2twLx9/COkMnL6gxhFJYPGaFFLAulXJPVL7yH31gFm0XcwdrTljMBGD1IHcIjtP
MY9FzaPFul5KycPnde+YviDxDN0pZKoEX750gcQDMURSFOuaYfmk+m3i0S7THeGd
vVJSFaFynC5lhP4w86sa0qTqEgKuDTMvbd4W+bs7KXlu9XInBEPjDsAUosSEaMCn
s1UkjgkmRwFBrIHxmk1Z+abXnmIaemCrGingt290ey8GjEUKA1xwxyuwDLaGfDSb
CYjlJLrsGip+uHPMzFSDcOwbYZstRa6Cc4RhtK6Ra1blXTol8UURn0S3xpbortYg
R9rmW8/Oj7dGwUZ3fudm5XXHVQ6+N9y0ShG+QohVPkFc5m0YGFugEKiKCq3XZJ/K
awhjqnmUvqpxYF4bKKtDjQx3Ya9poh8fWGn/o2AUYsnW3faP1Pzb1yxVOcJvpTtL
5JoA69CPOMeGQamX8aee9ce6mYHbYR95TeSBMlfTXmQpWCwROG1X75Gh/K2EuPeO
kcJ9i6NEGWlG2mkT9KDsK2bDEoDArLqikmJ/3CoqnblHpvTv+WviwLC+KSFlEdag
ceRBlNefwsKFvyZE2LfRSuovnlm6SysZ5RYX4+0pxJkDVAR5lCaEZLoJneVf0G+N
+bqbl3pGf84qegsgcohHOIizsIWdhokOjYrBYxccMhIor72fMr1nX03BJQ+mKXJb
IHh0DLbofq1cYBgLUUGWZWnoJZ+JaM1jjYKE68HgPYlUSWRxsWSH3ummuvLWx4ol
3lpjaDtom/VY0rXcbfVgRn7PJpMGFeWyE1TiDQJvG7AvimjEN7erVU5WpfzYCGd2
b2ipfBBnrreZGdEvnm+pJyWag6jWU+m3S9OgpeeT9BQS2z9Ct/gPz/x/WEXi26mK
5QECyHmUlYQ9CwS/ePSLLYnqrvnfNxnV6S0+sCTOhha5INdxJ001O+PZB4buMA93
miN2vsUc7JZqDQLPTai2Yn6rldZ1HO1dDtS9meClyR7rYcOikcw83qHpecRQcR6F
vE8M5pdRQwDmi6vWxPqMhu+yvu4RXaD6fOFewnPsLoHBAiqtJ3k3uHVL9DPYGj0E
NaWqggJw7sSMNt+pRQAYeOhfga2T5BRRlzZWiahi71Jao5qPWSbKSZxbt1hf17DE
87BxHFaO/wH7Fh4yh+cn8klD7SY1+C7cucKSUNH00cLctkiNMdzK2U3+bLFdojD9
W6VjJKl2fhh/AwgXAOv+/1gO0GNnj7zXxWJwWIIGUgPuripRVpfZL5KMBgoSd8yr
MTMMKiFOuk62ipgXWZKIXsUrwU0fl4ijrsfYvQWSS8ujfRVFUtBhB/1xab9HdwsZ
esrO4Qafc/1uaNgH9YUKogdSInRJdMAghOhRz3XFPLxW+KrdGHqHZA5yrnZqNSuB
WAwOzzdLJ3EMTpjvlNtkjzmXKwbSsSYmEXbAp6Rp3xPY9/QNXzQs8KKSA7nIJe6h
GXFIKTy9N5ggHj+IkPE/rdVC6/YKB5V6E5JSGG4ob6/IfSjxObgb/qBvr5tC/Tve
bMUvafZqCHPib73mOBPHCHydfzOgBcbql5D9KDRQ5fCa/uFHs65d47SYFdx9BbqW
EykGQRW+pPur/ykrBGNXAxYONWOiT58y2ZnIhMxdw/lZXdSG+QvSY/JoAHs1pSIs
ujFRZfDRzbZs1qlJGAQJoJLYRt+bfSEK4GmIrqQs3z3ljyXe+1SOuQfVFtfquGAT
hFy2niKKPYH6Pyj+4P02rh7c9WzImJIryzRhamTjH7zPl1ZLaXaKIXiY53TB1hxU
+LXg4G/VwdXjtb2v/40Lck3uvpsDPzY8OQFQbtJ8o5uIj7qiLDV30pqVDJOV0H11
SqiA6T/9yiSaXKzfH8ovSTLZaKQbrug8FuWRK8FXnDvy2YmT1yVDTrJlVmVPkAvY
hW8GLUzSUQ8fxaKRwSXQQNAATEJDZQoifL4CK88L1L8LoQ6n8YVUM8yPO9eXJVA2
G2aFmuBWzrX1qUHGRQw+V0qZzXoXZAkQnGB8rZbUuDi23BU+ZJJCiZ2hQ9qAABJU
LO8KoZ78f8vGWdHP6yQ786uZjTc/H5c+7TuExXrPc1XKaU4h0LfYgk9UYnbmIfc2
nN6aAsErSNcOoWf6IfX5N+ykaU9VsftyYNJ64AJO6QISrFiY+GMLc8tpeCVtm5H+
9mR4lyjoZZ52G4DfNSM1QUPy+cxoTpujYyAnM9TEBBXdnMb3p5a3cPHhTJKSp9CQ
uSmACRnqewtjlpGVNjKCDv0dKACBCGqV3MI+qAOP4QKBDwOF0MFTh2QnmjMtVVbU
5b6FKGtakHBNfTs828mSjSavZXzA77iftyjgRo8ltmEiO8Qkj1G6mYNJOBys/IU8
QNHmPxKx2Ty/oO2tBvfxwNNmR/Qwu+c8Nt/URB+ytTUkxJKc/dAKeR339zpejjRn
JE48yhBvQ14EM0sH0DqdS+KeTiyhri/vc6hsFhJqFq8k5cmlfNjnr7jNtkCpIEsZ
qa8desIWQBUcM+8oxM90lzbehVM7i7exur3E0U3oXj3wCwfqfjHtYDw3hXwrNldV
gukgT+vccdbPIRgzfVxy6cdHxv84ICCuVj0CBz4WlN54H9rRy6WqR5DzysYguu1k
qpodevVBg/GHI2TmbsP+ejRjQ6+oV2QP2zt5lL6+ww/ZPUjLDbg2tqHsP4Ls6LB7
i+Ktn1OlFoK5ZXG1HQKm87ZNgF00fBRHh4yvH3TwmEOviP6DS4rtqtpaLyt01Jak
b8yqoMo+xL1IR/8t6sZd8osyrDu1LoScLqi6vGL/orNjcGPXAOdxXygBpu+cf2Nl
utXQ1x7pfrkHDrhMgO4wkEjj5GFryDaXZBwQSqIqVckjfH6Un2ppQVFsAFOrQ69d
I8llVP3kCXwSUrlmjRzDIMsJvs9312S/nveo192KSVvOTQZT+Vc5XHqUU9skv8YE
8a18vIu9IEvwhw4RYGba6hRV+TSPfB5A70aAeox0S+xnfvmUwlwvJr/WOQ6L/dGk
Il3QtJrr0/RVXzxzV4mvfbE3vnYf7JkweYSmSYmc/nqDveqDjG2gxLtcUTp7fRe0
o9fvz+0xQw06H4Wlh8xsFa765TPc8jMio0kMGM6o1VGh0XPbdk+BZ9CHPeOirPup
bCKCIiDWDXFRz8i4hu9zkjAR7pgO2x1mpiJ7zMsjgNjIkV8Upta1v620M8PysU9H
l6HpVujlQeH3s7FBD4BWJ05TQvQWwHpWEqY2N0Wqw18HAxkuA1nYa97mel55iklJ
t1kCtQXn732Sst7A4uigdqJ4hqVHVliRhadUP0F9E6kXtUlYB0CO56pUVKocitmw
KCy41ScT32cWucOWNKhfFiCgfhGt12yvrDHuFqZ2ZKlb0PZe+Yz1okaHm/r4s6WZ
SB2pxZNlBbVjCV7w/aXMG7DJfV6EZspwB16h2xzQHUd2hiiIvstc2qIcPUaru2+f
DFQorKa6jWzGiSEA4WrEZjJWLDIvWwcLSTHM8ptRwGtwvkNhe8P8nOIped5cY5rf
c+sT3xxKytol89QTcsw5S30/tPeRVBKQ063WV4l/exbflPwGfQ7MzLTFTGVx38vl
dhxtTEgPAI+snRRHDUQTewdYHYAiP0xj1JkK4wZZBkt7AxK8vyS7bHpC86ndNNDh
Vwf38EW0HYEKoMxe6IAIDvLiZoOBFcamDDsmj43sX37SpuEaG74NoiK0ocJ8Cxqh
xzFo1RqvvCeeTtu5qjZ5LtRGrXwq3KsxLcpxw+xM8RH7hRjA3uOuoJa90fhQ76dG
Z82X95R6ElEOETEmQJV3OzcOm5U/zzwVKaRPAHz3pc68pf9im8eXEVgmYPvwUftC
fUzRMPmXPwck3nkppj6iOPrYWWWOuHtsupwpnlaCz0feeuGirnsll0Ij0p4vaxPe
bfwYE3dp/oEQ8zqOIgwME2Y3aW17Ik+qlM+C9UfBpitjq8KB8ulVDIZ0fLd9zBBV
0MEcXP5KVw1kQ3v3TImDhbvtzkAJF3QRXIF5kR/1eZu62PQ0FiOLc6wiiaPT+wz9
yDlhIgkDUoSzMYaXGkYb56moMtIVCWrZhuV2dyrU/v0/lwQsKlmhMpa0+Fa91XES
gKG8PWlxKqgGakKvpLyeQgGj3GyNNY0BgHhMA3NQR4miF6tUZc/aehPQgLwkG6Pw
1REoQIw4lwTVoCNYFBRCn3QCBr+y46SJt1XIR4IJi5L1ov5hp3Lp6FOUEEJrST00
nhMkwbsxPaDAuNUpU14waMu/2qCg1uDUs8bMAhIfqFRlOJpolHvFEaRUj0n2I/34
TdPiHOo/qbDceCJmuwfCXvfK1zgZd6ssq4L4WBPFjF0+V0XIACEv3NXRe7HWhOnN
rSBtP5hMn7zm6xVHKXhtQL/f9zU80G9MLt/fnVT35WqiFBp8kwZ5xMoyjvqFbu6N
bvjBAYSh0U7IttZR+6oAoxtO2ahZw1cksCQlqcK8FoVR4Ve29F8J22eazp4HPQSP
T5x2mvypxqpjqtaTMJGO/BjW9YlpxGL7qX7BH+blur/fN1ysL/n/LV4e0zYEHyxk
9EgjLP24WwuHfYqr3aX49IuXZ7U6L3uxwjYNdXGkQS8pL4Q/fhGUiMCaauu2ETkx
2RkzttfwHv5aJsmEEB6OadkOMs+srjMv70msqT8Zj1v79GgDfCncu3hGWDfU3OVu
OdcEYuGAI4VFPpoxFCxY7iN94Z1sj044eNVO3zLobsznJS9eieagLDWkWg1eqIjA
f8YIzDQAi9a391xtODTWWAwkUz5nuQUjKJJ/b60KXSM/Sx/kdmmDRDobw3WLbaRU
fEqPoE7XmprDFciv++yhs3n7l7QWLtM6+Du+ysjH+/cxh0K7KOfyuP4oK05Jf2Iw
j7MGMmy2C8Aw+h69UJWAQ0q4LYtqUeuob06et2Mdqo6n5wayGWudIx54Y90w5jq0
vh8xZGEPNAyWpCJOSDcd9xSRREr4h40af35MUB+WMorEowMHmpk/mllzCKQXmjju
D+gNosUGdBEWXZeR82e8qUXs+sKVhY5Sx7DuNti8ssJ1zZo2y7OBunCVIdzHcU19
Sc5USF6DkfMsWrOUDW5uNPhRP3B5gxkLLFEEoR0fGjNX7JpEut6UKNiz7h0aq8Ti
8dFmfN5Ptc24StaA02o8G5m8TAO2DypAio4leDrC30Echb1pOgpj3HTWGL21vnVf
GlXUXZ6U9HI2AmK+qujYbilnQxz7/eSStojG+SBvKzVcYuQjW6CfC6pbTBl3g2M3
2IuXvq0ZBf8YVtFJ2se+KczJT1LNBlEgBJoLy/DTAPziX8mSbT32CPg8aFDemg7u
gcpg7GrK9dZRi64R5HHiVWSfTWvBH6d5kpdY2Rd/eANX2tzU3Iz9Gu7wWK9J38eT
Crxc9/esRwiOXX5IEGptpHoEhASr8mNn4zkZnO6gTvudsY+YptGmZaz2YgscILCs
R0IRq0x/zE/XEA8E9lK24tHiTY+gKgTCWPM/Zuar3ZRQQw+q5i544YTNZ9LSdb8f
CbKC+6qWtubdMXCPY76cxHij8ZqTHEcJdWaSFNua7/iUzevg3HRk5tGuxwtmo0mj
ikQlcl0Img22DpeWid6HllXAlg75y8QVCnIXkSeLohOS6SF+H6yo5nXypVhRQ4a4
p04lO+7Bvf6rdwH7MKzF6LgUXZyo0WH2Ho/2tReve22qKjql1Zz4A5oeUECUj65X
WG+VPrgBpN2vzw+o9uENFcRraTQaXABv4qDXH4FyOD6c+9Z75U4QG0CJqEJsTjSh
1f+w+2KAsYGfIsESabDT6nOQuEt7DhC1A11vByfS1qYMQ/4u+e2PeEbwNnMuUZbt
RzLakkojlianrymVE3iVZDvd9lIqprXndV7njx0DTqYX8/p3iBPp253LU+5fsWTx
7eVv8nJKsUXzAZvaCHO3hii++HOJ+QKbNcQ45Igu3vS757csN6uZ0VPX7ENJhAeS
MOI22IoGRFkn6ubKxuChuUszhi37xjdIiw6F0vWvq4HDcLEa0HevlCVmsHnus9RA
krPZRrx8v3gOJFNzPB1Bwiu8WqKtDTSij3ySag6EQCB19oiaMfOKgK4lJLGLd/k9
cktNX66aAds7/xYyxO1wDxPRevYJJNetW0UJtrDtno8uvl1B+u1FXGIUU9JsduUq
EoBnbuPmFOTiELpHepPFZ4G6bD6GuGFsRZLk18jjuLX1u3fGWp8yVjbrSI7cRdTN
CVAgyYjZ7U9joSpM/wVTHk+Quo8PIpijhrTgUFhZdWyBFWLCvQDjWRwGvbo/jmYP
Db0Cg4tKzHglb0Z0GnAi/rKBz4HB/+/jpaaJ9jWT6hGDpnYgSkCYZoIOTn4LbkOa
oXgIyLUe1gPwaJChxaMoepmlkB2FFrVLk4+5eZjJjgSdmk9ysD5eCrPUnR1MObEv
Lo/F4Z0WxIESIcjHcpe75e559odIEkgJ+R8lnnatOZE4wiVyMqFIstSukGEyb4fZ
j2U7vN04ZKb5WOmTMNIQ4Nr/WPQLe4C0ePaI6/wmW+SBNLqWqkiNJOodQFQoJq4w
F4EKZojboiw5yrRge/MTd1QQUDCSjoTfJe4IBlUq/sfm57yIf+Yx+udv7cfHpYQ4
FKsKu1jB9RkpREo8k+wFxcjkh8OeyKNZ//NuGTJm+9oMJDg4Ono3eqwnBJM4gtcA
EA0V4Awd1g923Y4+0zXPUHhh6acYNI8wV6FswPBt/K8aCB7y3aFycVO2SwZ2XPU2
ylsbrOeSDH/4MVlMH2V3cKUIysOJQwwxyxGhSJhV6Y15+WKrEcVzZTvPKgb4y7O8
7QpKAZs1xImHWTTROB7I7ELi9OdxTVzVRdWqxPBjj6hfC9fGZRyTF0GmpLkVXBfo
AF/2V+NzliGKTFZ1jT+Mw8mO1wTJjK6Q+Bo4gGAeOuJw0zpDIujgiLSaAZmQX8JV
IGFcQiEkXKOUjI8KjwU6m1reUXafrxIWE6U8U7bQS2t2zWx/t7rwC5g+WrQo1VT7
l2zkZTcHm8kqrTMQNCWKeNyN58IjjmHAYsdIQUBxMQ1lIexK/yfutGmZSu/fQzly
XNWRdXSUi/upwrCLyt1iW3iwksYnPkr4ZnU8u3+/anFqi6iOM3nqfFBL+fJxAbm8
VmdSIV7GNVHbkf3E9CHksNt+SR7fFXC+k6IEkLZpmxIPP+L72vA1aaZkshMGuZXr
NxzfZ324aGMAVZwSJOe820+M0eCG3Wv9D9gLJEiV7cpzv+0pSYqlgi+NSc8MQ3ve
rq82LPLPl0SwV5zbXa2u1OxzCAv3RJ+iYUJsNS/bbmFm7t9TSS89t4LcYL/2JdWP
UWN9eqLgqOKjMF+Eu4M19uTMMWeEB6sf4OHBaqYS0w1CctZYFxHNuwljthFNr3nf
qKqlpM7YYRtf7YOli0kpm+tambe2JoJc3ppC9WndmFO0nUPBIheulqx2ddOwCXgF
KEIcMmkf5e9UWLmyt8oY7cmpTVDqCyO3lPhNea42foRXL+riME6oT3BavmljEXFm
rH/KSDceMbDb85ixtEcVm19EkSp+T3LR0A5rp6DCdj9r0DmhMk1rEGwNcx9vWbQ1
RNnhZ9w0cV7VzbRLs+L35Bkog9lQzkvnHRlQfG+cYg1TuJMEBpckM232iQ8aJhtH
SMpDEMIviChHYSdPW7G0d43BgnbiYHQT2SxOxy9TCFbmw9QTzn7aLJ9VFe9IHR4P
6AsPJw6iVz1fZi7JSnCp20Rkh2ZBIvPDNAcs4KiRE7L0gM4HiYAuMVttUmDs0l1Z
fQalPAqe+aQbbsLEyKVz+jGTr7445tgcNFuuVNQe6m7C5R7OMqPCpFrlL2Tel9OL
QslYXaquGnSVrXErK/aH3if+/UjLELhFhRAEpilR16qKLSu8dJ2fyFOgE24ibsR9
e/455D75cMt7vyYAROQBH58ZHkW8+ZpweR+CdrsoRCIfdixhnv1jaZOJqS/Lh1wt
nkolo9UayzG4oRTIukjaawA7x21Wyc3k8VqIKdVZieWRawOX/mDeMN9DRgWOcoS0
IV1fQgklG0L0YzCYZNOjwthErab361UPTgOwUY/BicPmjsimJs4XrQdKzpMIX+cz
xII48xGQAHddv++dBXZs2fcO2Xzuh+9UUEm+FwrT6nMDjj43ggUrfGonhtR4aOnO
Mf73ljhGtaQ85v7bPmJDxYJcYefUVJbnjSY4C+KH77TtYKgrzRG0TzNQ8YhSVC0j
gYX2Xw1U6xtiDuFN6GKDZJ8sGRtPz7BIYQ5xsPlRKbNdsrXRR09CzURb0Vg65lVQ
OauSa71PBjdKYIC+Ke2ZtQZSJchLI3vhZAaMuuAfVlS0EWhyzo4inR3wL/AQMaaJ
hx2lha4N+nS84uoQrljbrcCUpqlqiKa+zLMQqSdc6fVG4uHsz+uD5aPTJym0bQxw
jQX/RHBL6xj8H3A1vD0r9XGWZLSE3yeN04c7YNxNz+L5IwW9PhCeCvcZcR7tiXIS
iZtzQAc/X0Ff7IKehuLubAlU8elv7tBJwogJvX4puaHB5XVsqqlSkSZi/xecJvKe
9mP2TDqKiMlb96VfEO0hCXGRBb6/f7eo/modTXBdoQj2/Ym05sRVYlI22l6zY9tt
fZKO+q4FIOjwhSYkfexMlpQUShhUagpe8hIjROAP69NFvUl4Oy7X53doWSS4S3Yz
NK5zJGUnaChx0E5Ikrz0ObkQVmObVzSQfGZXRSWzA2adFR+UWkFGxAJ/toOOpS7+
mr3MY8HHRBN1MZfFpiDITWUpOlVv0jSU88lADtXPdEwxfSyX/uRHtb7OfaAefDrO
nImw32dv/0c3bTiEScyUJs4UQ8kxgU2VHME4+Q+VQUEkpJBri1lo5EiWpxOMsUNM
xIWwAsBViMDPBNCuq2Z8qMGqLO1AP7HUL0rQ9pqhtJCtn70rq5Y6Ztw1fnj/ksJN
v98aZYHpLVAoUdDCdsA3XtADiMRqVbKj1650UevaGSLWC3tRCaz5XzOxeWnF5Btd
9LXiWsM2K1zmgZg04Wc/dS26tgiy0lsL1u6vTTnHuBFmHCHeNz97Lk4/1qGRUul8
/HStLMCdZp7Wb64kpkVNVL2F4JRr1ITEAe8AytgYgzMAhNsJiVTxi7ySU+H7xs8e
ZsJb4jMEq3MGD3H8eLPul3OKkEh/R2mOdb2qoX0YR/rHxZ8snPUErd5Kroyj62Xj
EH4DMorRhH2Rxb23k0O+IdhfVH2t0LNpSYWM01AB2L2y+x8kMPgwmFK/wE1C7WKz
8w4NaZkRcwEBFf9aPxPHWNgWqLdHGl/TcNNb88wCTVcvX15GLXy68z9BtFke5PNH
/4H0mks9AmXxUc5/SFnG/Ky1lMwa1dOtD6JOiy7yB4HByfxu1SV+EtOY8V2ScofT
grkICgFLX5hRzL3cgUWLxgU0vzUlPoE98CSoIu7T/ZBIqeMIX9H6sh8sNyHgS/z4
+uWGBk58mSc0hXdyPQ8c9RKyr0NCL1H/f9lZqfp1opiVWk2oMUjAP+dAgn4CNDh9
zWh4yKb/ZjKEGdgFwfUHjE7HuNzxC9HrvPU7D/bT05k+P1rwqG8HBhuBfmMhBXfL
ctqNH/1Yh39bzx3Jx6lrdZSD5lTZZh6UZpol7PoxNxcWy0shIRPBWvu/dZHKEagQ
df4vBY0MF4Zks4MROAowao/dqz7Mapz+bEIATpOdpgfJ01LTLiJC/Ns4QmjuL1W4
UZY8sVLYqtAFbQIhc2Lnzh1Jocigq9jF1RlIZoabeJjip+uF06/slhV3Cfz+bfzz
FD1f946UFchz8uf1mxOj7Ljmcrlvju0qpGRmF9h/zE9RQbN6FrG9xNRMcnL2Hrks
rDD2ERcx9mDcc6vZdwXZQDrO8LNz0d1AHwchlf1vRFkMLxrMx/8cxq5YUWIuTqPR
oMJuKnAJwJXyf3sbL1Q+1sePb+fI1pEjwWRMzuE0bMAyXuwzz5ejRJd5FK7HXXmg
T4cgz8zLK+r8KZ1Fa+uhTDQsBlGkWLGqWNO0TxgtCleYTmo6byF7RCb1maV7c3Rf
b4NKEXpdqcCFKi4sGpdVUyh7yNEVuCorCzdkW+lTokDrWLeaEoeQ4A9E3VjlHVG9
pLSIBriG6jUE4kshap6AJ/AWKqFGSYo1G+7MV7W8JqYZoPXM9D8pJbsjEGL1dP8O
h+ntRNiJtCqo7rf2HELWTWcjill6IJQbMcBZ+SToRHk1nRJ7qmYL1ka6DIZPd67X
WQmPiF8xQyWqVFdITcaZJnPjAZNfsGs9IyslDvR06AFeI14zWX776j0YBbyV+reC
Hew11b7ovWfMKvSgEnvpTyJVNIcLMw6wd71N/QMQVHJM5uqNTzAsh87UyESTJd+d
97dVYFLeAt6945+XT4WM2Ed9wqF3vkkHlQ3jEHMweDhySHIsnTPeu5iZw912gUif
XNJ3tQ4SdMKs34GEkuL7F2F3yMrRO/uELWYiBPbdCobu1RcbcTfDy3pnzZVD2mgj
pZWp/XRzWxlkSIZOBxPgCwrSwAk9uOb67b+4EtQ2NTh/irp8JcopWTDauFjBebZB
/87rcGmjRTVSLQwNbe7xZUbfASGwZJ3vFbI2fV3cozXtwoEynYtYeCgKIDzS2JLO
o/k735JMKux0jVjlxSYbojXIxGk72La3geRirv1orifiyVD2m9hQFtBN92MNV4Kh
bz4pdur3emH6fYUTnWV7PDSgn6/wtyaaqK3BVLIHmzsBjpOyAS1wfqTxnK7fbgid
58Lw0C9zDjZrjVvquwIVwSvKRrutnJYFHg8w2fpaOhkIkTCEu0IjlXAjYMV/vU2y
meeqy0PW3aCpg4z6uh4+aIAa9Si9pU9QF1ZxMMIxor/hfP/zrDbloIEr5uWMdPIj
nSyd2yuiIRhrjh2C3iWFnK4Z9WcDytwE8Q1k42s8N3GE184+Tp0RAGNOxuCiyjSt
9UTNJEgN3ipeFMRe9NtnbcIXo/jIB2tNJ9ytiJu7MVk3HHp4jQBP63VpVIUsAbFZ
DLEmkbacn/T2BoiJtmU3HLR+CKILdY5W8oCtOtOKqTXnE7TWo/OAplP7cIGta/VS
kw4ygo8SjPROgq9cv1qlody8LIf4EAJS9LAWaEAB9Q6gcNk6aWvL4KlFsgM9YvGz
AotolYBYxX8OuBV82gZLHp0/wnA1lLPd3P7FwYkMYhXjPryXKdT4EQLrU5P9IAG3
pZSYkDoHkuRVxei6zXBWecPSA3O4nKRV6Q0wbtVW9p1DyPypgGdCNUKGBTRlVfuw
uE0wkLECXnw+ODm0jtGNE+KwbMuSdq+YnXpjKQxLWbIai6brdrMLaQ8hss2qRMM+
r5SQPrOHjaOOW7rPsrspcQLftH2Mh+WYiB+furcVjiNREg4vNaOrzqzxGV1F/jFd
a1tLFLYmBgQfNPVgFXtr0mG83SeX63l52jm2Ya8sKfJUTlVDmqsKQyuzT+OrGmMP
6yQOzLYPyGcZO76GszvMBq+gdOgA1Zqo2BPcixKJ4w1uoLsQ0VzemyN0WRHorXDH
+LFDBzAStOpMtg8VyvqYCQbnqIq2ggx5RNXIf/M2VSuIlVlhI0C9BrZb7p31G1W9
mwPqky+6EB+8ZuHw31XRZpGs7m02G0BpOusjJPcOP5Ht2fBrmzU7kwcLX8xTAItB
KoqIh+1xbf53eg+RGTOfDzPnDprJtt+ih0sq5p4++Z2Yx5Z0059Vxtj2SLPq92IL
6zyyThTmmOSRsfKJzX9F/nFRcJLfnfuBXZhyIMr8/i5HMkkIuFR5GWv8TFWu3pYU
oZdVZGYXO5BgV3jse3RhaG4/0UmNwf8UhNShAVTWbsrxV1pkZgeskvB/fZl3tRnx
0qYBTpQLj6/ZYnx5sf0TSCHx26/JgFj7lEpBHvAtkuw0dfqwmcTYgbln3fDoy0Ga
8mNP7K4aK329tFxawWWxAZWq/5oQWAza7Us6arHA7V0Omb2LFCg5xz91d0PvuqqF
k4FXKPsrHszaAT9UyKoALzC7xL2qTl+QqiL0BRbmFvWFg/lmFKLJQQRR+GQVq7zd
EfTc6pkXL7igYWkbEkey9R6B0/qj5ocwRM+IYdxsFTkELMhDLq24a4no9szr9cJ6
KUPCm5Xuz2RADBlQ70XoSA6fsR0X8IIj96b9mDhvh010CB/fTCingf1hfaNCb5dt
9U45PrpUyMygP4eAPaGq8BUUyEzAYDgyU3SG8gE2uWQrO9yFhvRAcXhWFyYedgD0
o9wJROtPSJfI/v5tuDAfLtpGEMRk6yfOP2rrIrusPYuYfePOO5bAU+Ns+Cnv1mCw
8G3nnCp/AZqvxnXWsp5Kx4xjOm5kzQHochq01R5qM/H68EAFcx2D7I0UUWpBwISz
kXspqKLoHA6uEZWWxXA13PfA8LIdhljnORs7/mcFXNjqDSJbQTFZnyGNPbJ/cNzl
9tFMFxnzTg6nJ0yD3X+YlvqwOixvctQnygMpwUbqGRceAJjcQMY6qCiGF4ww/l+Q
NQYYyrnR06CQkzqZikFz5xfu6Iboy2PR8XTpf05qZL0an+mIO1HvYJAgW/bad7TP
Ppq7UNtg4J1mgwU0Opxp8Q+P3VugYRDXZeRe6c6iIrfinRFpmDV6kGWHtw4L5L2p
QyGleJl1VHbT/qesTmpTVRePvSqneeJqpra/TaeyV2BBWbbTmG7Ydw9B0J6oSGYH
GTpIQr+0w1StdgbzUQIlAyo1O7tpyv3Jmq70ZNqKpm8A3zAItv2i0s+4LpI+KK/q
SxE55gX+wy24TE0GkH7bw8R3Xqz6eksi2yKMzRDPexSeOkhVKOXmbKakyhE3hz/N
fAEq5pAL3/17MKr+dcHo/9fdxiDAmo31aAumg7hxcrsWvM/N5PuTVjZp94ZPQKxW
OFQkNiysMnETwKwh0B4rRQKv6y8+Hxhbuh+fqWbxwLvaASUkk2NZ7BwfuYH8c8Ga
GNlUp8OE1QOq/VuLHs8UEHW5YUbGNl2HP+D4HXGGJqDpkDvfJuznqrS5dseD5oRc
fvvJHzttTHpPvbRAIa182GVPhISJ9ARqKhdU+X8Yd2lGrvI0XlF1I6BZziPLmHe/
I8ifMRRFjQ+kkWWf/a3zLUW+JqmuszrXfaRzISYMAgup8RuDcC4apm0xExRPTqsz
XKCN5vJrkxwBcc9prscd8BvCeZXgiZ5NlySnOfzBRXCs93gUl4MFCk0CIw49X5FA
2D0m3hlqxi2EwqVDzRevFE9qDrDB10lrDkZEzDWxanfI5twcL57dThovNwUgADRl
gnLbIaFNYWrKOTFWR0i/qKr4OjDLovicHdELl9VFTnoD4sKnT84klp1egoF4iStl
f0Hm8cpfTvm4IZaPGcIaPt1fFTK1JDfAZsV1xL1qlE/URglBxYjkAYcgo7q+fV9R
uZYbBkBVsNF3tA0Ts3mOH/hacnrHDUsSN9WTm/M42ppmKCz9QQOory/zPd2jJJPO
GRhTk7BzKdYtk4hcxvQQp68CZwfEKSS07zAxuh1R33zJmcaqCcHfRUDZMckizEqm
6H02X0TI9qXK3UWUJ7UTr61R6tvZKVvfDl6fjKPPexNe+k9HekboHYkxLtH01vbd
s5cb/KMZzpLviP12QosPQ8dY4gKPBOxPwlGTJf8em7iNUNTrbcyp3DbOT6lRfP13
BNAK9R9T+By5zRaQ1vt/a+iJsuWkLcQ/eN0SzJ7ntr9t/xwwNmgBPMcjMYZl+xsL
vv+Mlf6Cii6nrlG81UV4BsXrXI9UQX6LIYA3H8E6ZREB8zBj6axqdjJ6ewLJAkN1
CLoZMJ4sm+YxIcGMCN6Icv8Ar6ZEuJzWZBs9TaEKFDxTTmq5rK5bMNb/sNh1P6Pt
Rcuoa8VLfsDZjl1+d4gLyOo77ViqwF9JF3fZrqBDAIXmGP4WCYV0uJhI/lq3tort
Bmm/BaQlL0TRQ5MwoACiO1HAI5+KPKRAG0/ZKhZaeNfKY5CX9G6Swk6jZYlPkQmJ
Lf6Y1Xn1eoABVML6/osLY9RDV+pMjC01tJqn5yNDKF3P+w1fsNcGmuu9sK4RKTH4
zJ7DNXTkxuXz/Tss0jfW8LlyOLlWaRNR5jzwB/LRWUpJbiqEQLFsy30wGHkb7UmX
sJrw2LWQaE/BGyeIul9NdvqCTaQ9RXQ7A+pKL0T7Z9X4RcnBi1xPJM6+7Gs95fqs
YENxVLwfW+xkeBe7nItFNgDtfdAo+Zl9RXWLuRXjIAHVaKb/J1sBAP/jfXqwIMWL
NHNzChVlU4O0SFMRpOg7iFR6t8sWHjed2dFXmu7XKzm5B8GDUUbgkQwqWG8bTP0T
hfcfb+QsdPA+O43x/eoMB+G1Sns77DoE9fQOQq3RzufNXr6mA/FOWQsAnCE6pHga
SnaVb+xRShnw53keS/uadbBKWecIOLUNL1lgq6/sLJzzYBhQ5bh8/rEB+DQuc+JD
75I1/C/nmLp+lPQDjjeOQ/W1G0xMPUYvnMS8rlkxh0UY8MoyZIjNwSnNhgQW35Ty
tvocmwXKRBzXlJXJ/E0Sr5giXIheugjZRtu5rmyWfQ10ioiEmH9+OvGzjJYv+LkJ
VX9nqNOFUKws2gYK57FwlgkhNSNfXHC1jMs+Yk4wp8g5jigNCZ9P5X2vcO9ijgi/
N9ORhMuRPb0VEeqF/YBtvkLsr+zoOqIT3OLUTuKTbXG1bH+HKKtB82D+1Lfrgg55
44ppWNrsnj57OEhom+b2iK9aEgP04qrG/DLFer0jG+r7dVHRNn2TN5lnQzVhtyrv
J0iFwY7cb/TvRgB7sKI4cOSCFb46YjKjn5XpkFyOfW9z4oi4dytQRwY1HeinUiVW
UpC0kImahhNbknUZKI6bC0IUdkyQVknNqqSxSju08RyXTLW+WhLPWWshuZkJe2t/
uDvFGrSH96jy+Ucd/fBsO4IOAzcIyMcCjKXELkOwtBso7xyIAA1MeCiYSC9aKcRV
K3/lrBHXcZPmtpUqzEegW7niC0Pk19/ubvhDCuM3ArR0As/t4N7+ghl0aLAxLE07
kYcGNmKjPKwR3o2YcNtwDdPMD0RZAWbm95Zf7jnLyOGIPzeVJKbnvn4YHmqPd3Zf
GmN5vHZaXSfMwQ4wM1qAUeefGSMMR/BDlVMdx36lU0dUXhmu5xNRvnnOzHH1bXix
QTi1zk81yCZau6IlAxXw9UpC/q5WBYsDOzlSxPSRc27S4dQSHLuTx/X6ubMaCsY4
yFWxaTZ9eL9YgKAFQzc0VSBegch4k8xLEivhAYSxt8HIhszypDxtGUQJMw89fDO2
dbTltLBtFdCaLINhDpqC7oV2RwMdAMRuJHKXIUH/nQ6SyKWEVy/yPhuZb88QrKyM
B1lw4sSp4d61Z0G1eC8ZQQU++MqGUucYsZBDBBwduidpaLI2FPk8bXzefjCwCRmb
RSnH/0BpJ/jDdXNbOHdrdXlEaTqqzDWcr+7NddJ2MxOvmn0BI9jlQAQS3//jGb+v
wz/dJ2ghK2mlJqj4daNzawM9H3u1A7rtx041rSarmNadjRAi3WLLh99+d3YRiQEm
DcecmVzarfVCxyZF+whxHBS/y/Jac+wqkGq3HIRV/6gTFXySqX0qDgmjzGh7jwiH
MJsRH7OfDKD6L62UF/zwXjSHnT3wCagSUpL2L7OWbVUUY+OsLeNj3ru0LdP3FcQK
pAQaxioq7IQrgTg6zucs6KP7xsCxBbE0TF2mwz1bQ01QmhQ5Y0LZbADh8gFhRvAF
N0M0mFPgMMYmbw//dSY6qWUEoBb7ezEVci636O1IYMa7v4iZDslJBTHCRYFyDqi8
9bCY5r2fuVSk2QI9Xeendm/ChWojoAzlM6Jy+j+aHbEYTnoMy8f+x4lBRu2gd9Ir
UwZsOzumqjk05JobYiOYctz50iJTYcdcI/zeXTazjbVlLdXCBw57R1avxkRB7FBO
eo2UAqOin1D8NqcyfT916iASnweJRZqAvht2Fqvej2xHEfkuabSIDdoXRZlaRr/a
APprfT/WVezIur0ouY4BO2hgRx9/x73LqI45ABXmQdpaULfSz6h7hhWq3nk0XbGX
ZgzSHhgoRepijUkPSZGdvSrYFO9A2WB6uDxim9o5Q4q1N4z8dr0Ib+s6fIQ6Y2LY
5ghZrbpWSeVsxA2YbzQR/GA18tU2MIB5g3gzjaV7zPKXzksb0FIlfor/D01WjwUO
BfypLt/QVFB4tF90o2U1ScUD9dPOJfi0gmoZMQkDD5QucEnSV1ndPUcUH/BSofP7
P5YcWkXpxTj/uFS510LIVmjJ7R9P917CR0sP/J/sZORCHIa2CC7GTZzB2LRMZ8/J
NNW1ZPwmIDfJP1Md0CZGfnpNaLAzCFjCM4U80/Be/lvvyHMj6zqP2taw/sZ1djby
UKMOjiogxx5aEZGTUOtJ04CJXar/rZUNOh7oedqyn6QvKi/+XCiG/btGowKSiUlB
0Pq6aOwYPKoUC7QvT95brNviIvS58Uxb1pQgG4Pjm06NKnQW1nGSra3OXuigllou
R2dFcr8G114UkkLWY2K6tcMCnsBlZchRKcqP8zN3D6xVczUfMIhlCHmi5K2N8+qW
6fXUB4HRUqC3rL7HGB1MBdJxS3BNUHJ6BIfsGsbKdomzrCDEkInYlic3+HTTc8W9
NsP7NG2YzwQlEAq6/v/pJjSLWoU7DIcuSGwuny6jvi9bmlae6MHP85wnXd+vzJLa
aIuzsGw8+n3WWqvJKmAo5k7sY7p6zWQLbHhWMQZyWbOpyOxtiXaRFtaoLHZma7DZ
ZU3Kl8h3xA0nze7PTiPcdyjDGPdSnv45FwgbC0aIRD6bBuXq5iZWXMIpV3Fg/lZw
j7lzh6PzndnAI69HneaEP3rXnUe0zOxOwXviL7npae/IHqMYQ9PPA8hgMZNIfb59
lCH9Vzi/YbxvlRV73eL/6lN4YpFYcKAmny7I619ufpHp9frv8ZhwgymeDM/JdnlZ
/Ao2cW35dqRlDDClrUZI7mBwlDB2ICzAAJD1bkrT/AsEFeq2C5pvKxzV6rkqvV5b
el9AFAjhuVl4yDKl3GS9eiMyjjgIk9fxt0LiPY2WMSCcXXnODui4exGV6mcdJ5M6
rrJ3a4CadRN1nM15g1YRsiR3374UE5z5mV8ZMpIJ4WHAdmRAh8RV+ft2SZlbvLbz
xg26mo3pTlM8voCdinTvoptk+SrfX6p05A0mhA4DDvk/PfXelsas47Ov6Gtm47XI
30R4qZPjrv1sCC0zMoUcsvrSH+gkdSch0XYYoI3SZ0/UTk8epbFe8fJUnCMZMCLg
oV8LYGTL1skfpqu612d5chw7/hHkH+0DuMb+R3JUNUasOecnuG0QlhfiPB4oIqFm
m7IFZYoRGC+/Dez5JsOUjHJFo0sml8OvYQ7S3/vm2GYyJqfHM+7oE9dUSPtiuzGJ
vzK2XhMoYQwGxAul8xmwPcDMva/LbVSloU20GTvCi2WeJjKT7qHyJVlNMOeMr7T9
BUEE2+ysf3kyzcTtYfVU3GORCVGF2Li4vmP2XqbaRIPgWgrCv1LBquqQQoNobqZ+
IgIxCyzMvMYsaGEVz7tgygmMjD2wGuU4M7H1K1NQEBH0eMseKmxVyI/W0BE9aRAU
RNCpCFLrHVdJbPn1t9O7kegEvlxESbzcWQbdsu5fn/JkUz2JD3qBeZdiEN8GleTj
Y8UF5sTYt1WYtIdNjMAQW8/s1NP4ON2nCIhXOYY8oWFw1AuuL2ohsLsmc3bWdcxu
pV3tz+r5OxnmLFskAwTdGf7DrytBltPH94Meb3NktBh8T7d61SYZ89fku7okNrKB
zsBcWORA13TpntfyaX441CY7bwJHZhigReIn7JeP/x+Zjh56DQ+I2//lIC4jWzaa
+YL0hukN0cB5C1SmQ4HYncjsz9L10QlkpI4xScSw8fr1/bp6RfkJjUeizkxl+KzI
FEC6y+vFeR5RynTrz8bUxlL4/QtJ+KgsKco2r2OvDHdLs/BHL1164XPhTQ2d0njy
oXo9fDX5eA3RP5g29XyoCmHbApDYpqbdZhevgFpiq7p72YJkAuV0eAbveWQ2y6IX
gozPwJIPNLngm7vB9wjm16wCdTXCH84o2rUeUAuto/bb2ZaBbdknm9vUJlYTFYDo
oAfSXC+/FSIqoQmnai9PkTHiebJO1tcerSTrhrcDTNkELWaVcOi9/QyiMHoZVNDs
J4tl87ujDzuEGXsKBZBp5NfCoUz7RDWvWwlNBek3u9geQMnj1WnkGRYKT6ohzuAc
VBMY8NS04SVL8RKEp0LaZ2EQpWH/3VtFg892pqnU8FJOWpgpQb4S3YMk9j85ZGOo
+wGCA2FeYdt+YJE3tL+V8eu66GI5SN1bYhZcbM7ACXHPaUWCNzmSC+BPwWXpgXkI
BwfGpkZaumZAMDMaTQ9MS+bMSzn2pR857B55YHvfdBwuVrt328fsv7oBkGumTS5v
PXeB7XW1oUGuOrdfW9vA3Tmbz35E7ePk42dnXMAWqb/eJo30HGRDd+5lUaraEn4n
9PQAlWyiQMobxzeOijpuPk0HJEsEMJwv0vgdz7jwOTUiRIebg1LC8d6UZ8SJmFnU
jyTznUc3CQF/Xn8xy19oTYlwh+LpeXLQKJ4Vo4OhQzFzyTr83520Ruvjp6RFJuJu
oahceT2snHksOtlTmi9LTGoZBtaW1SD4jPvwb7q1uBS9lgouVv9nlUotzNGnPW/3
JNlq+/mqU9RkVRAgGdyfU6KU7QK6i1tjNCI9YN335AI9NfeNOKeyvTkgDxZKu23S
1WaXeJWwLWohqcICI4uccw/kjIPCYusUzZ44pf5OGCwJ3BFX/BHh/HGd+SLRmILi
O/ldOXvxZuFD1NUx48FTciviQ0el9qFNa3dT2zI0FPntxLy1igfdkdWsW2MC9cfq
+lsscdVkgTuzvi8V1k6elBOTqTIogyu0AfDksGdtlnanW+E2iFq7b76ZSQEF2Air
xZ1wxLkFh3jj0BJV6k4nstusjQvD9fGsnezamuaG2trEBdbyfKKXXuM/iepaTCrH
s2UpcohJSmsNpV0EZbFZlFMvmRPA3UYPxBg34uidO26ZPSBh2KbPxV5CGICufaF+
qAnb8LWJhvN6hW83+YeL8v4vwMbc0qGu0/IqPCddPf9p0dUO8GUH2Ka0fnNoz1CQ
c0owEVDPiyqS6uL7Yqlr8r+YaH1HORKqUTif0Uh6Oe3pyW0CfK+SsHrUweVQBXLk
H3NqohiGzOfw5nt1fAQ0YFdF4JJT9hU+JCRtCLy5qkg/5mDFW5YKa4GsyHXAdy6H
1FrVADuwU0casyCKa6i4fPVpraSz/X+nHCGf7avr6z/UlIlIYdHHdJ/hFfLbP7FJ
daqiaq1IUJ7mEe1XG5duxd2lMOjmFhajZBeaioB+dQ2hoPXAfI1+0eaJjNAltnJl
MrLQ3JAsJt0Qge/4dRx1tk13vGMPzIOaDa5wao+gLoiffKFVlC4Dqrx/wZS7Tkic
oeZVhg2gsJ+bPrVlKU8Iratu/SFfMcq/nuFpjXfUCYE4nFEcs15UCU4x1VSM9bdq
0sMiQpQJB7K6cibQv9xcWWnJVuD/pIKS1fkRgMIOWJaMCS1N6hQypxoIkOy4tXAW
QhjhMfV+tKvOdm4d1MS2RWVIobGSoUfolmzY5Szr1W7+GJmLnj8vxxUypOpSyamu
oxTigUhkmncn3zTOJJBaL5NM4HXPfuZbf3IZDVRb4JQ/VNbQtR9ldJAFew+cVZo9
WgJRbv72CTMDkDjKjQ2zzGtOLQBaUnKd8Qz7Pe0eRi+f4KIwzGXo7ravCk14ZSfi
7x0q0kGDTEk56vuit9qWBHllUKDua5gd/PLeCcm2jOP5tP6Bynqfl/WL634ntBdZ
LjtV1yT2SBZebibvHr48QcqRI9h6fwYLWGtl/6skEjHP1j/V7+X84P2s0GQjP/n8
f/9jxjzJv1o8X+BBX0F2plidEpmUuV/lgYzG1vc7VFik/GLJ0QmTn2TC8eTr33sv
xxNlf/hI2QS8EQ6821URs/IF/lzM1Wbs5JS81kWFnF8UK18eQL43pjbE/Cx1oFY7
O0Fmr909B4OoXFQn82UK6rptYfO8AZWW0IiWajXijUgFnLntXB2QOa4uMfU/SAf9
UZEw6v1MLEkZtYzHt2ySM8KyQWWugH4SqIZdOKid7w+5qYa4urwtxZS8953ANdLS
1kSjblGDI8OqDGmkfFCO035B/bu4twYJdaJzwo8zAAm5/JBzGNvWzaP/wQAtmlQc
lKxWHY0O0v4fA2bzaetRajo0uF2m051uq0DAdxvfcuZJ6mzpeD785AHAtN3FfBED
OiF2ZLKa5AeSS+QVbM9Gtub0x7gkFkaPjUX+6jR1QQQZVVJjNeA0vV4df0C6ifBF
DrJzkxLt5ZIbuomlau8OM1L5L/B9ZvQLZvJQCKqJCdRZzMFAU8GjZ8SSCwx+ZU3h
9oxL/ldOWM6CloQlGl4Qeb3GY9v3JuqSB7j6eSK4b5FAH8wIPuWYI+sbTR8/X+aC
KB2sybfw3HVpBfcSpx9hTt2ME6Vynk1yTRDNH1Ol8QHH85uLoynQlNUbAlMH7Omk
TbkvBTZVrIoGD9kxw2x6XB5BzGSO1maHBZCmUDW1TYngFK3xvP47L3bcoh6IUpej
EXCPZuAs+dvnGjhlN3FtJoNxbwDwH8Ylst2Fz4ymkl1zJaaQVp3dVvWLY7nMrLQP
LVCy6gKKM0aPquYMDC8D3uTxKzTiL81WZ0OcQKyjcVeV5yQnVGd+jj/zSebvz2+4
95QR2fzhv7Y/Pk8tDsdy5gvnfE8Bx/JCAAx+Vb2PydorW1qRKe0L8WwcrJKM0ME7
C5uCybsjQEFVl3k2c8jeuiu1sOpFsgeEZnOddwJbmn19saTwQzM/+l7QsKavL4GL
2ArSf2GZpCfO+5eoQ76Xkv132aIX3EZnG8ZlvTiUSEotoEtSnZMmXL56WQZQSmDi
ESozg7ya5daCNpOh81ug5OqCapijzNbplgtNkO8mf3PaAnBrwzVqCuSlculG5ImA
cm0ipS0XXigEXVF9rFvvxs08ef0oYayro+jNymYKKFWb8fmUzcc3S3JpjXfvA9hL
C0u00iVDK5z0khK1UFgc2ZJUWNQ4Qvj1QlL/Cl+7hEMsGD1DQs6isNxti8Y4+AVc
vL3zjIV5wq0u68b7Q3P/IhUBdc0qdfmePRqspMEf+cwXrlFwLzgx3yMIJk+/NEGP
47NlxMap57Hjp8y4ZUncTsfJm4hz2gtU6MzeQtwcW3hR7I1sARNSS29ASQ+hnF0n
aFuDZ/ocG1qYsTNwfhYl/IMdLL8pvn9Y9Oi30QwVmLF1DIHpbnY1zFgK2UVyyF4v
G+O7T+SmpsCmgCKdopCf+utrLgyu3vbw4qz9Yu3ZqwQPYL8vNaQ8/JrCJwZG0LPF
2pr0G1E7w9+LmWl+UJRdZSzndhZcvknTdS6OA+IKuyrp9bqGBgClEZJ+JMukOcAa
ujBZ6fj+ji/26rwNs7qAnT8lzVhkb/+yyB2j1+0EVJ5Nz4oQvQll+xfMMJJOWzZT
OqPS9KaJh3/QWsdERX9sVwA5+R4ahY4v1kRLxgN/1tdkq/6M1Xg8UPMlP1sGwl8S
K3/Dlx9+EnU70EjmBc7fk4f2Xi9lTixAUiNdqRvcyKfC7ma4zUUL/AtWs0IjPrWr
aPJkacnWOAN/YGbPSXm28tR/acmVQQH7wrLKrSOxpl+bl4v2WoOU4O9S91f3KG7O
g8HvKwzmx48pxzFG/lhCTztwBWUe8/TEN0VlmFxYaC2H55410JWNno6j162uzDgm
FvoIh5gTf/mkWVroHY4mD5waabbKh99GFK7N4rb2CVBL+xuSe9pI8PagEcqtBtGR
oTiEvDsyhZbM2IC/U3c7ncZg606fkxhZtsmyrQXNa/RhvxkKe4E5X2DDc/c0z0R9
kEeRdgnPL2HdCBKDL30PH3+j8uWep6C1qwjPmuUP7NyXkEFwuAHm3FvQeee4S1m4
H84JwqnTmoVEce7QnFZ4G9wqsG8OQA4OJBXi/+RfYUXks8mUW+AKgn0a3lAKC8Qd
czY+kUf4fs6jksMCQB5hHkuGqH5AZ76DJk1qAtH9iT4vsOAVt+Z248sxBlPfGYUs
xtI1Wm3wbVbBDpL7lcA9H0O1fmV1vbT5tK4oOELlGTfA9NSLLt1Xa9fSAD41gpd0
8kI9Xp0lXNUsSxZ4o2DHbQ35MbEGZfiumnRgf8csDVDwpWUNa6/HwohmKFmPWuTB
WHJq6v1xOkQVGeEw3kdgGkOYMqvMcKg/0q7B9XxGehtJIaNZbbtXcS4CX+DGKlPa
Fm7SbLZoaG/d45F6bwLhcN9Rh30fmpOswCfQtqsiwVy+BZgUArlcTGP8tfjqSEPy
2+HdqrdscD2pcu5MIHDivzhiHEGM9zVJVaoIWtgu+TLawyG150hGdwcV8KETEv/y
07qJRrhPwIEw0c2MWMEmvH38+6TDyRcDRhhuesfZ0/6Ed4P4avTxKorGcY/WQd4N
DaZnoFf7NfAXetJfVXKWv4Rr9Hha7gmX7vVlXViF9nA0/1H7lEOzFLQhR9C+zS8Q
JgYSji8Wuoq2gMxZ+ihw0ICxNgtIBt1qgTTJUF3P2KgwBqG5rKoUM+fJ4J78dLlz
iCZLRXla2IpkTruwVqT9Jwm3CgNo6wrcK+Rz6Eh2kW4=
`protect END_PROTECTED
